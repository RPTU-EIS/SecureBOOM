module upec_miter (
  input clock,
  input reset,
  input [63:0] data,
  input [63:0] secret1,
  input [63:0] secret2,
  input commit_index
  );

  parameter PROTECTED_ADDR = 32'h8abcde00;
  parameter SECRET_TAG = PROTECTED_ADDR[31:12];

  wire         auto_intsink_in_sync_0_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_int_in_xing_in_2_sync_0_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_int_in_xing_in_1_sync_0_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_int_in_xing_in_0_sync_0_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_int_in_xing_in_0_sync_1_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_a_ready_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_a_valid_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_a_bits_opcode_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_a_bits_param_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [3:0]  auto_tl_master_xing_out_a_bits_size_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_a_bits_source_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [31:0] auto_tl_master_xing_out_a_bits_address_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [7:0]  auto_tl_master_xing_out_a_bits_mask_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [63:0] auto_tl_master_xing_out_a_bits_data_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_a_bits_corrupt_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_b_ready_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_b_valid_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [1:0]  auto_tl_master_xing_out_b_bits_param_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [31:0] auto_tl_master_xing_out_b_bits_address_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_c_ready_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_c_valid_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_c_bits_opcode_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_c_bits_param_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [3:0]  auto_tl_master_xing_out_c_bits_size_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_c_bits_source_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [31:0] auto_tl_master_xing_out_c_bits_address_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [63:0] auto_tl_master_xing_out_c_bits_data_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_c_bits_corrupt_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_d_ready_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_d_valid_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [2:0]  auto_tl_master_xing_out_d_bits_opcode_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [1:0]  auto_tl_master_xing_out_d_bits_param_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [3:0]  auto_tl_master_xing_out_d_bits_size_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [2:0]  auto_tl_master_xing_out_d_bits_source_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [2:0]  auto_tl_master_xing_out_d_bits_sink_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_d_bits_denied_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [63:0] auto_tl_master_xing_out_d_bits_data_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_d_bits_corrupt_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_e_ready_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_e_valid_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_e_bits_sink_1; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]


  wire         auto_intsink_in_sync_0_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_int_in_xing_in_2_sync_0_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_int_in_xing_in_1_sync_0_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_int_in_xing_in_0_sync_0_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_int_in_xing_in_0_sync_1_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_a_ready_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_a_valid_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_a_bits_opcode_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_a_bits_param_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [3:0]  auto_tl_master_xing_out_a_bits_size_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_a_bits_source_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [31:0] auto_tl_master_xing_out_a_bits_address_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [7:0]  auto_tl_master_xing_out_a_bits_mask_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [63:0] auto_tl_master_xing_out_a_bits_data_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_a_bits_corrupt_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_b_ready_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_b_valid_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [1:0]  auto_tl_master_xing_out_b_bits_param_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [31:0] auto_tl_master_xing_out_b_bits_address_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_c_ready_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_c_valid_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_c_bits_opcode_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_c_bits_param_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [3:0]  auto_tl_master_xing_out_c_bits_size_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_c_bits_source_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [31:0] auto_tl_master_xing_out_c_bits_address_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [63:0] auto_tl_master_xing_out_c_bits_data_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_c_bits_corrupt_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_d_ready_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_d_valid_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [2:0]  auto_tl_master_xing_out_d_bits_opcode_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [1:0]  auto_tl_master_xing_out_d_bits_param_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [3:0]  auto_tl_master_xing_out_d_bits_size_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [2:0]  auto_tl_master_xing_out_d_bits_source_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [2:0]  auto_tl_master_xing_out_d_bits_sink_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_d_bits_denied_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire  [63:0] auto_tl_master_xing_out_d_bits_data_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire         auto_tl_master_xing_out_d_bits_corrupt_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_e_ready_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire        auto_tl_master_xing_out_e_valid_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
  wire [2:0]  auto_tl_master_xing_out_e_bits_sink_2; // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]



  assign auto_int_in_xing_in_2_sync_0_1 = 1'b0;
	assign auto_int_in_xing_in_1_sync_0_1 = 1'b0;
	assign auto_int_in_xing_in_0_sync_0_1 = 1'b0;
	assign auto_int_in_xing_in_0_sync_1_1 = 1'b0;
  assign auto_intsink_in_sync_0_1 = 1'b0;


  assign auto_int_in_xing_in_2_sync_0_2 = 1'b0;
	assign auto_int_in_xing_in_1_sync_0_2 = 1'b0;
	assign auto_int_in_xing_in_0_sync_0_2 = 1'b0;
	assign auto_int_in_xing_in_0_sync_1_2 = 1'b0;
  assign auto_intsink_in_sync_0_2 = 1'b0;


//Instantiation of SoC1
  BoomTile soc1(
		.clock(clock), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410017.4]
		.reset(reset), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410018.4]
		.auto_intsink_in_sync_0(auto_intsink_in_sync_0_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_int_in_xing_in_2_sync_0(auto_int_in_xing_in_2_sync_0_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_int_in_xing_in_1_sync_0(auto_int_in_xing_in_1_sync_0_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_int_in_xing_in_0_sync_0(auto_int_in_xing_in_0_sync_0_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_int_in_xing_in_0_sync_1(auto_int_in_xing_in_0_sync_1_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_ready(auto_tl_master_xing_out_a_ready_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_valid(auto_tl_master_xing_out_a_valid_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_opcode(auto_tl_master_xing_out_a_bits_opcode_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_param(auto_tl_master_xing_out_a_bits_param_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_size(auto_tl_master_xing_out_a_bits_size_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_source(auto_tl_master_xing_out_a_bits_source_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_address(auto_tl_master_xing_out_a_bits_address_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_mask(auto_tl_master_xing_out_a_bits_mask_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_data(auto_tl_master_xing_out_a_bits_data_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_corrupt(auto_tl_master_xing_out_a_bits_corrupt_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_b_ready(auto_tl_master_xing_out_b_ready_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_b_valid(auto_tl_master_xing_out_b_valid_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_b_bits_param(auto_tl_master_xing_out_b_bits_param_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_b_bits_address(auto_tl_master_xing_out_b_bits_address_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_ready(auto_tl_master_xing_out_c_ready_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_valid(auto_tl_master_xing_out_c_valid_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_opcode(auto_tl_master_xing_out_c_bits_opcode_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_param(auto_tl_master_xing_out_c_bits_param_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_size(auto_tl_master_xing_out_c_bits_size_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_source(auto_tl_master_xing_out_c_bits_source_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_address(auto_tl_master_xing_out_c_bits_address_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_data(auto_tl_master_xing_out_c_bits_data_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_corrupt(auto_tl_master_xing_out_c_bits_corrupt_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_ready(auto_tl_master_xing_out_d_ready_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_valid(auto_tl_master_xing_out_d_valid_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_opcode(auto_tl_master_xing_out_d_bits_opcode_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_param(auto_tl_master_xing_out_d_bits_param_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_size(auto_tl_master_xing_out_d_bits_size_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_source(auto_tl_master_xing_out_d_bits_source_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_sink(auto_tl_master_xing_out_d_bits_sink_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_denied(auto_tl_master_xing_out_d_bits_denied_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_data(auto_tl_master_xing_out_d_bits_data_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_corrupt(auto_tl_master_xing_out_d_bits_corrupt_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_e_valid(auto_tl_master_xing_out_e_valid_1), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_e_bits_sink(auto_tl_master_xing_out_e_bits_sink_1) // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
	);

  //Instantiation of Memory1
  TLMem #(.PROTECTED_ADDR(PROTECTED_ADDR)) mem1(
    .clock(clock),
    .reset(reset),
    .data(data),
    .secret(secret1),
    .auto_sync_xing_out_a_ready(auto_tl_master_xing_out_a_ready_1),
    .auto_sync_xing_out_a_valid(auto_tl_master_xing_out_a_valid_1),
    .auto_sync_xing_out_a_bits_opcode(auto_tl_master_xing_out_a_bits_opcode_1),
    .auto_sync_xing_out_a_bits_param(auto_tl_master_xing_out_a_bits_param_1),
    .auto_sync_xing_out_a_bits_size(auto_tl_master_xing_out_a_bits_size_1),
    .auto_sync_xing_out_a_bits_source(auto_tl_master_xing_out_a_bits_source_1),
    .auto_sync_xing_out_a_bits_address(auto_tl_master_xing_out_a_bits_address_1),
    .auto_sync_xing_out_a_bits_mask(auto_tl_master_xing_out_a_bits_mask_1),
    .auto_sync_xing_out_a_bits_data(auto_tl_master_xing_out_a_bits_data_1),
    .auto_sync_xing_out_b_ready(auto_tl_master_xing_out_b_ready_1),
    .auto_sync_xing_out_b_valid(auto_tl_master_xing_out_b_valid_1),
    .auto_sync_xing_out_b_bits_param(auto_tl_master_xing_out_b_bits_param_1),
    .auto_sync_xing_out_b_bits_address(auto_tl_master_xing_out_b_bits_address_1),
    .auto_sync_xing_out_c_ready(auto_tl_master_xing_out_c_ready_1),
    .auto_sync_xing_out_c_valid(auto_tl_master_xing_out_c_valid_1),
    .auto_sync_xing_out_c_bits_opcode(auto_tl_master_xing_out_c_bits_opcode_1),
    .auto_sync_xing_out_c_bits_size(auto_tl_master_xing_out_c_bits_size_1),
    .auto_sync_xing_out_c_bits_source(auto_tl_master_xing_out_c_bits_source_1),
    .auto_sync_xing_out_c_bits_address(auto_tl_master_xing_out_c_bits_address_1),
    .auto_sync_xing_out_c_bits_data(auto_tl_master_xing_out_c_bits_data_1),
    .auto_sync_xing_out_d_ready(auto_tl_master_xing_out_d_ready_1),
    .auto_sync_xing_out_d_valid(auto_tl_master_xing_out_d_valid_1),
    .auto_sync_xing_out_d_bits_opcode(auto_tl_master_xing_out_d_bits_opcode_1),
    .auto_sync_xing_out_d_bits_param(auto_tl_master_xing_out_d_bits_param_1),
    .auto_sync_xing_out_d_bits_size(auto_tl_master_xing_out_d_bits_size_1),
    .auto_sync_xing_out_d_bits_source(auto_tl_master_xing_out_d_bits_source_1),
    .auto_sync_xing_out_d_bits_sink(auto_tl_master_xing_out_d_bits_sink_1),
    .auto_sync_xing_out_d_bits_data(auto_tl_master_xing_out_d_bits_data_1),
    .auto_sync_xing_out_d_bits_error(auto_tl_master_xing_out_d_bits_denied_1),
    .auto_sync_xing_out_e_ready(auto_tl_master_xing_out_e_ready_1),
    .auto_sync_xing_out_e_valid(auto_tl_master_xing_out_e_valid_1),
    .auto_sync_xing_out_e_bits_sink(auto_tl_master_xing_out_e_bits_sink_1)
  );

	assign auto_tl_master_xing_out_d_bits_corrupt_1 = auto_tl_master_xing_out_d_bits_denied_1;

  //Instantiation of SoC2
  BoomTile soc2(
		.clock(clock), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410017.4]
		.reset(reset), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410018.4]
		.auto_intsink_in_sync_0(auto_intsink_in_sync_0_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_int_in_xing_in_2_sync_0(auto_int_in_xing_in_2_sync_0_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_int_in_xing_in_1_sync_0(auto_int_in_xing_in_1_sync_0_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_int_in_xing_in_0_sync_0(auto_int_in_xing_in_0_sync_0_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_int_in_xing_in_0_sync_1(auto_int_in_xing_in_0_sync_1_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_ready(auto_tl_master_xing_out_a_ready_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_valid(auto_tl_master_xing_out_a_valid_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_opcode(auto_tl_master_xing_out_a_bits_opcode_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_param(auto_tl_master_xing_out_a_bits_param_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_size(auto_tl_master_xing_out_a_bits_size_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_source(auto_tl_master_xing_out_a_bits_source_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_address(auto_tl_master_xing_out_a_bits_address_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_mask(auto_tl_master_xing_out_a_bits_mask_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_data(auto_tl_master_xing_out_a_bits_data_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_a_bits_corrupt(auto_tl_master_xing_out_a_bits_corrupt_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_b_ready(auto_tl_master_xing_out_b_ready_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_b_valid(auto_tl_master_xing_out_b_valid_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_b_bits_param(auto_tl_master_xing_out_b_bits_param_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_b_bits_address(auto_tl_master_xing_out_b_bits_address_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_ready(auto_tl_master_xing_out_c_ready_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_valid(auto_tl_master_xing_out_c_valid_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_opcode(auto_tl_master_xing_out_c_bits_opcode_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_param(auto_tl_master_xing_out_c_bits_param_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_size(auto_tl_master_xing_out_c_bits_size_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_source(auto_tl_master_xing_out_c_bits_source_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_address(auto_tl_master_xing_out_c_bits_address_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_data(auto_tl_master_xing_out_c_bits_data_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_c_bits_corrupt(auto_tl_master_xing_out_c_bits_corrupt_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_ready(auto_tl_master_xing_out_d_ready_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_valid(auto_tl_master_xing_out_d_valid_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_opcode(auto_tl_master_xing_out_d_bits_opcode_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_param(auto_tl_master_xing_out_d_bits_param_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_size(auto_tl_master_xing_out_d_bits_size_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_source(auto_tl_master_xing_out_d_bits_source_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_sink(auto_tl_master_xing_out_d_bits_sink_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_denied(auto_tl_master_xing_out_d_bits_denied_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_data(auto_tl_master_xing_out_d_bits_data_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_d_bits_corrupt(auto_tl_master_xing_out_d_bits_corrupt_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_e_valid(auto_tl_master_xing_out_e_valid_2), // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
		.auto_tl_master_xing_out_e_bits_sink(auto_tl_master_xing_out_e_bits_sink_2) // @[:chipyard.TestHarness.MediumBoomConfig.fir@410019.4]
	);

  //Instantiation of Memory2
  TLMem #(.PROTECTED_ADDR(PROTECTED_ADDR)) mem2(
    .clock(clock),
    .reset(reset),
    .data(data),
    .secret(secret2),
    .auto_sync_xing_out_a_ready(auto_tl_master_xing_out_a_ready_2),
    .auto_sync_xing_out_a_valid(auto_tl_master_xing_out_a_valid_2),
    .auto_sync_xing_out_a_bits_opcode(auto_tl_master_xing_out_a_bits_opcode_2),
    .auto_sync_xing_out_a_bits_param(auto_tl_master_xing_out_a_bits_param_2),
    .auto_sync_xing_out_a_bits_size(auto_tl_master_xing_out_a_bits_size_2),
    .auto_sync_xing_out_a_bits_source(auto_tl_master_xing_out_a_bits_source_2),
    .auto_sync_xing_out_a_bits_address(auto_tl_master_xing_out_a_bits_address_2),
    .auto_sync_xing_out_a_bits_mask(auto_tl_master_xing_out_a_bits_mask_2),
    .auto_sync_xing_out_a_bits_data(auto_tl_master_xing_out_a_bits_data_2),
    .auto_sync_xing_out_b_ready(auto_tl_master_xing_out_b_ready_2),
    .auto_sync_xing_out_b_valid(auto_tl_master_xing_out_b_valid_2),
    .auto_sync_xing_out_b_bits_param(auto_tl_master_xing_out_b_bits_param_2),
    .auto_sync_xing_out_b_bits_address(auto_tl_master_xing_out_b_bits_address_2),
    .auto_sync_xing_out_c_ready(auto_tl_master_xing_out_c_ready_2),
    .auto_sync_xing_out_c_valid(auto_tl_master_xing_out_c_valid_2),
    .auto_sync_xing_out_c_bits_opcode(auto_tl_master_xing_out_c_bits_opcode_2),
    .auto_sync_xing_out_c_bits_size(auto_tl_master_xing_out_c_bits_size_2),
    .auto_sync_xing_out_c_bits_source(auto_tl_master_xing_out_c_bits_source_2),
    .auto_sync_xing_out_c_bits_address(auto_tl_master_xing_out_c_bits_address_2),
    .auto_sync_xing_out_c_bits_data(auto_tl_master_xing_out_c_bits_data_2),
    .auto_sync_xing_out_d_ready(auto_tl_master_xing_out_d_ready_2),
    .auto_sync_xing_out_d_valid(auto_tl_master_xing_out_d_valid_2),
    .auto_sync_xing_out_d_bits_opcode(auto_tl_master_xing_out_d_bits_opcode_2),
    .auto_sync_xing_out_d_bits_param(auto_tl_master_xing_out_d_bits_param_2),
    .auto_sync_xing_out_d_bits_size(auto_tl_master_xing_out_d_bits_size_2),
    .auto_sync_xing_out_d_bits_source(auto_tl_master_xing_out_d_bits_source_2),
    .auto_sync_xing_out_d_bits_sink(auto_tl_master_xing_out_d_bits_sink_2),
    .auto_sync_xing_out_d_bits_data(auto_tl_master_xing_out_d_bits_data_2),
    .auto_sync_xing_out_d_bits_error(auto_tl_master_xing_out_d_bits_denied_2),
    .auto_sync_xing_out_e_ready(auto_tl_master_xing_out_e_ready_2),
    .auto_sync_xing_out_e_valid(auto_tl_master_xing_out_e_valid_2),
    .auto_sync_xing_out_e_bits_sink(auto_tl_master_xing_out_e_bits_sink_2)
  );

	assign auto_tl_master_xing_out_d_bits_corrupt_2 = auto_tl_master_xing_out_d_bits_denied_2;

//*************MicroEquivalence**************//
// Some info on ROB: it always commit a full row (two uop at a time), uop in
// the same row does not necessarily have the same br tag (mask)
//
// Is pnr (point of no return) important? pnr should always be after head and
// before root_id
//
//For which of them do we need to check both instances?

//Function that returns if the given ID in the ROB is a branch instruction
	function automatic isSpi; // should check for both br and j and jal and jalr?
		input [5:0] id;
		begin
			isSpi = ( (id == 6'b000000) ? soc1.core.rob.rob_uop__0_is_br   : 1'b1 ) &&
							( (id == 6'b000001) ? soc1.core.rob.rob_uop_1_0_is_br   : 1'b1 ) &&
							( (id == 6'b000010) ? soc1.core.rob.rob_uop__1_is_br   : 1'b1 ) &&
							( (id == 6'b000011) ? soc1.core.rob.rob_uop_1_1_is_br   : 1'b1 ) &&
							( (id == 6'b000100) ? soc1.core.rob.rob_uop__2_is_br   : 1'b1 ) &&
							( (id == 6'b000101) ? soc1.core.rob.rob_uop_1_2_is_br   : 1'b1 ) &&
							( (id == 6'b000110) ? soc1.core.rob.rob_uop__3_is_br   : 1'b1 ) &&
							( (id == 6'b000111) ? soc1.core.rob.rob_uop_1_3_is_br   : 1'b1 ) &&
							( (id == 6'b001000) ? soc1.core.rob.rob_uop__4_is_br   : 1'b1 ) &&
							( (id == 6'b001001) ? soc1.core.rob.rob_uop_1_4_is_br   : 1'b1 ) &&
							( (id == 6'b001010) ? soc1.core.rob.rob_uop__5_is_br   : 1'b1 ) &&
							( (id == 6'b001011) ? soc1.core.rob.rob_uop_1_5_is_br   : 1'b1 ) &&
							( (id == 6'b001100) ? soc1.core.rob.rob_uop__6_is_br   : 1'b1 ) &&
							( (id == 6'b001101) ? soc1.core.rob.rob_uop_1_6_is_br   : 1'b1 ) &&
							( (id == 6'b001110) ? soc1.core.rob.rob_uop__7_is_br   : 1'b1 ) &&
							( (id == 6'b001111) ? soc1.core.rob.rob_uop_1_7_is_br   : 1'b1 ) &&
							( (id == 6'b010000) ? soc1.core.rob.rob_uop__8_is_br   : 1'b1 ) &&
							( (id == 6'b010001) ? soc1.core.rob.rob_uop_1_8_is_br   : 1'b1 ) &&
							( (id == 6'b010010) ? soc1.core.rob.rob_uop__9_is_br   : 1'b1 ) &&
							( (id == 6'b010011) ? soc1.core.rob.rob_uop_1_9_is_br   : 1'b1 ) &&
							( (id == 6'b010100) ? soc1.core.rob.rob_uop__10_is_br   : 1'b1 ) &&
							( (id == 6'b010101) ? soc1.core.rob.rob_uop_1_10_is_br   : 1'b1 ) &&
							( (id == 6'b010110) ? soc1.core.rob.rob_uop__11_is_br   : 1'b1 ) &&
							( (id == 6'b010111) ? soc1.core.rob.rob_uop_1_11_is_br   : 1'b1 ) &&
							( (id == 6'b011000) ? soc1.core.rob.rob_uop__12_is_br   : 1'b1 ) &&
							( (id == 6'b011001) ? soc1.core.rob.rob_uop_1_12_is_br   : 1'b1 ) &&
							( (id == 6'b011010) ? soc1.core.rob.rob_uop__13_is_br   : 1'b1 ) &&
							( (id == 6'b011011) ? soc1.core.rob.rob_uop_1_13_is_br   : 1'b1 ) &&
							( (id == 6'b011100) ? soc1.core.rob.rob_uop__14_is_br   : 1'b1 ) &&
							( (id == 6'b011101) ? soc1.core.rob.rob_uop_1_14_is_br   : 1'b1 ) &&
							( (id == 6'b011110) ? soc1.core.rob.rob_uop__15_is_br   : 1'b1 ) &&
							( (id == 6'b011111) ? soc1.core.rob.rob_uop_1_15_is_br   : 1'b1 ) &&
							( (id == 6'b100000) ? soc1.core.rob.rob_uop__16_is_br   : 1'b1 ) &&
							( (id == 6'b100001) ? soc1.core.rob.rob_uop_1_16_is_br   : 1'b1 ) &&
							( (id == 6'b100010) ? soc1.core.rob.rob_uop__17_is_br   : 1'b1 ) &&
							( (id == 6'b100011) ? soc1.core.rob.rob_uop_1_17_is_br   : 1'b1 ) &&
							( (id == 6'b100100) ? soc1.core.rob.rob_uop__18_is_br   : 1'b1 ) &&
							( (id == 6'b100101) ? soc1.core.rob.rob_uop_1_18_is_br   : 1'b1 ) &&
							( (id == 6'b100110) ? soc1.core.rob.rob_uop__19_is_br   : 1'b1 ) &&
							( (id == 6'b100111) ? soc1.core.rob.rob_uop_1_19_is_br   : 1'b1 ) &&
							( (id == 6'b101000) ? soc1.core.rob.rob_uop__20_is_br   : 1'b1 ) &&
							( (id == 6'b101001) ? soc1.core.rob.rob_uop_1_20_is_br   : 1'b1 ) &&
							( (id == 6'b101010) ? soc1.core.rob.rob_uop__21_is_br   : 1'b1 ) &&
							( (id == 6'b101011) ? soc1.core.rob.rob_uop_1_21_is_br   : 1'b1 ) &&
							( (id == 6'b101100) ? soc1.core.rob.rob_uop__22_is_br   : 1'b1 ) &&
							( (id == 6'b101101) ? soc1.core.rob.rob_uop_1_22_is_br   : 1'b1 ) &&
							( (id == 6'b101110) ? soc1.core.rob.rob_uop__23_is_br   : 1'b1 ) &&
							( (id == 6'b101111) ? soc1.core.rob.rob_uop_1_23_is_br   : 1'b1 ) &&
							( (id == 6'b110000) ? soc1.core.rob.rob_uop__24_is_br   : 1'b1 ) &&
							( (id == 6'b110001) ? soc1.core.rob.rob_uop_1_24_is_br   : 1'b1 ) &&
							( (id == 6'b110010) ? soc1.core.rob.rob_uop__25_is_br   : 1'b1 ) &&
							( (id == 6'b110011) ? soc1.core.rob.rob_uop_1_25_is_br   : 1'b1 ) &&
							( (id == 6'b110100) ? soc1.core.rob.rob_uop__26_is_br   : 1'b1 ) &&
							( (id == 6'b110101) ? soc1.core.rob.rob_uop_1_26_is_br   : 1'b1 ) &&
							( (id == 6'b110110) ? soc1.core.rob.rob_uop__27_is_br   : 1'b1 ) &&
							( (id == 6'b110111) ? soc1.core.rob.rob_uop_1_27_is_br   : 1'b1 ) &&
							( (id == 6'b111000) ? soc1.core.rob.rob_uop__28_is_br   : 1'b1 ) &&
							( (id == 6'b111001) ? soc1.core.rob.rob_uop_1_28_is_br   : 1'b1 ) &&
							( (id == 6'b111010) ? soc1.core.rob.rob_uop__29_is_br   : 1'b1 ) &&
							( (id == 6'b111011) ? soc1.core.rob.rob_uop_1_29_is_br   : 1'b1 ) &&
							( (id == 6'b111100) ? soc1.core.rob.rob_uop__30_is_br   : 1'b1 ) &&
							( (id == 6'b111101) ? soc1.core.rob.rob_uop_1_30_is_br   : 1'b1 ) &&
							( (id == 6'b111110) ? soc1.core.rob.rob_uop__31_is_br   : 1'b1 ) &&
							( (id == 6'b111111) ? soc1.core.rob.rob_uop_1_31_is_br   : 1'b1 ) &&
// soc2
							( (id == 6'b000000) ? soc2.core.rob.rob_uop__0_is_br   : 1'b1 ) &&
							( (id == 6'b000001) ? soc2.core.rob.rob_uop_1_0_is_br   : 1'b1 ) &&
							( (id == 6'b000010) ? soc2.core.rob.rob_uop__1_is_br   : 1'b1 ) &&
							( (id == 6'b000011) ? soc2.core.rob.rob_uop_1_1_is_br   : 1'b1 ) &&
							( (id == 6'b000100) ? soc2.core.rob.rob_uop__2_is_br   : 1'b1 ) &&
							( (id == 6'b000101) ? soc2.core.rob.rob_uop_1_2_is_br   : 1'b1 ) &&
							( (id == 6'b000110) ? soc2.core.rob.rob_uop__3_is_br   : 1'b1 ) &&
							( (id == 6'b000111) ? soc2.core.rob.rob_uop_1_3_is_br   : 1'b1 ) &&
							( (id == 6'b001000) ? soc2.core.rob.rob_uop__4_is_br   : 1'b1 ) &&
							( (id == 6'b001001) ? soc2.core.rob.rob_uop_1_4_is_br   : 1'b1 ) &&
							( (id == 6'b001010) ? soc2.core.rob.rob_uop__5_is_br   : 1'b1 ) &&
							( (id == 6'b001011) ? soc2.core.rob.rob_uop_1_5_is_br   : 1'b1 ) &&
							( (id == 6'b001100) ? soc2.core.rob.rob_uop__6_is_br   : 1'b1 ) &&
							( (id == 6'b001101) ? soc2.core.rob.rob_uop_1_6_is_br   : 1'b1 ) &&
							( (id == 6'b001110) ? soc2.core.rob.rob_uop__7_is_br   : 1'b1 ) &&
							( (id == 6'b001111) ? soc2.core.rob.rob_uop_1_7_is_br   : 1'b1 ) &&
							( (id == 6'b010000) ? soc2.core.rob.rob_uop__8_is_br   : 1'b1 ) &&
							( (id == 6'b010001) ? soc2.core.rob.rob_uop_1_8_is_br   : 1'b1 ) &&
							( (id == 6'b010010) ? soc2.core.rob.rob_uop__9_is_br   : 1'b1 ) &&
							( (id == 6'b010011) ? soc2.core.rob.rob_uop_1_9_is_br   : 1'b1 ) &&
							( (id == 6'b010100) ? soc2.core.rob.rob_uop__10_is_br   : 1'b1 ) &&
							( (id == 6'b010101) ? soc2.core.rob.rob_uop_1_10_is_br   : 1'b1 ) &&
							( (id == 6'b010110) ? soc2.core.rob.rob_uop__11_is_br   : 1'b1 ) &&
							( (id == 6'b010111) ? soc2.core.rob.rob_uop_1_11_is_br   : 1'b1 ) &&
							( (id == 6'b011000) ? soc2.core.rob.rob_uop__12_is_br   : 1'b1 ) &&
							( (id == 6'b011001) ? soc2.core.rob.rob_uop_1_12_is_br   : 1'b1 ) &&
							( (id == 6'b011010) ? soc2.core.rob.rob_uop__13_is_br   : 1'b1 ) &&
							( (id == 6'b011011) ? soc2.core.rob.rob_uop_1_13_is_br   : 1'b1 ) &&
							( (id == 6'b011100) ? soc2.core.rob.rob_uop__14_is_br   : 1'b1 ) &&
							( (id == 6'b011101) ? soc2.core.rob.rob_uop_1_14_is_br   : 1'b1 ) &&
							( (id == 6'b011110) ? soc2.core.rob.rob_uop__15_is_br   : 1'b1 ) &&
							( (id == 6'b011111) ? soc2.core.rob.rob_uop_1_15_is_br   : 1'b1 ) &&
							( (id == 6'b100000) ? soc2.core.rob.rob_uop__16_is_br   : 1'b1 ) &&
							( (id == 6'b100001) ? soc2.core.rob.rob_uop_1_16_is_br   : 1'b1 ) &&
							( (id == 6'b100010) ? soc2.core.rob.rob_uop__17_is_br   : 1'b1 ) &&
							( (id == 6'b100011) ? soc2.core.rob.rob_uop_1_17_is_br   : 1'b1 ) &&
							( (id == 6'b100100) ? soc2.core.rob.rob_uop__18_is_br   : 1'b1 ) &&
							( (id == 6'b100101) ? soc2.core.rob.rob_uop_1_18_is_br   : 1'b1 ) &&
							( (id == 6'b100110) ? soc2.core.rob.rob_uop__19_is_br   : 1'b1 ) &&
							( (id == 6'b100111) ? soc2.core.rob.rob_uop_1_19_is_br   : 1'b1 ) &&
							( (id == 6'b101000) ? soc2.core.rob.rob_uop__20_is_br   : 1'b1 ) &&
							( (id == 6'b101001) ? soc2.core.rob.rob_uop_1_20_is_br   : 1'b1 ) &&
							( (id == 6'b101010) ? soc2.core.rob.rob_uop__21_is_br   : 1'b1 ) &&
							( (id == 6'b101011) ? soc2.core.rob.rob_uop_1_21_is_br   : 1'b1 ) &&
							( (id == 6'b101100) ? soc2.core.rob.rob_uop__22_is_br   : 1'b1 ) &&
							( (id == 6'b101101) ? soc2.core.rob.rob_uop_1_22_is_br   : 1'b1 ) &&
							( (id == 6'b101110) ? soc2.core.rob.rob_uop__23_is_br   : 1'b1 ) &&
							( (id == 6'b101111) ? soc2.core.rob.rob_uop_1_23_is_br   : 1'b1 ) &&
							( (id == 6'b110000) ? soc2.core.rob.rob_uop__24_is_br   : 1'b1 ) &&
							( (id == 6'b110001) ? soc2.core.rob.rob_uop_1_24_is_br   : 1'b1 ) &&
							( (id == 6'b110010) ? soc2.core.rob.rob_uop__25_is_br   : 1'b1 ) &&
							( (id == 6'b110011) ? soc2.core.rob.rob_uop_1_25_is_br   : 1'b1 ) &&
							( (id == 6'b110100) ? soc2.core.rob.rob_uop__26_is_br   : 1'b1 ) &&
							( (id == 6'b110101) ? soc2.core.rob.rob_uop_1_26_is_br   : 1'b1 ) &&
							( (id == 6'b110110) ? soc2.core.rob.rob_uop__27_is_br   : 1'b1 ) &&
							( (id == 6'b110111) ? soc2.core.rob.rob_uop_1_27_is_br   : 1'b1 ) &&
							( (id == 6'b111000) ? soc2.core.rob.rob_uop__28_is_br   : 1'b1 ) &&
							( (id == 6'b111001) ? soc2.core.rob.rob_uop_1_28_is_br   : 1'b1 ) &&
							( (id == 6'b111010) ? soc2.core.rob.rob_uop__29_is_br   : 1'b1 ) &&
							( (id == 6'b111011) ? soc2.core.rob.rob_uop_1_29_is_br   : 1'b1 ) &&
							( (id == 6'b111100) ? soc2.core.rob.rob_uop__30_is_br   : 1'b1 ) &&
							( (id == 6'b111101) ? soc2.core.rob.rob_uop_1_30_is_br   : 1'b1 ) &&
							( (id == 6'b111110) ? soc2.core.rob.rob_uop__31_is_br   : 1'b1 ) &&
							( (id == 6'b111111) ? soc2.core.rob.rob_uop_1_31_is_br   : 1'b1 );
		end
	endfunction

//Function that returns if the given ID in the ROB in SoC1 has its busy bit set
	function automatic isPending_1;
		input [5:0] id;
		begin
			isPending_1 = ( (id == 6'b000000) ? soc1.core.rob.rob_bsy__0 : 1'b1 ) &&
										( (id == 6'b000001) ? soc1.core.rob.rob_bsy_1_0 : 1'b1 ) &&
										( (id == 6'b000010) ? soc1.core.rob.rob_bsy__1 : 1'b1 ) &&
										( (id == 6'b000011) ? soc1.core.rob.rob_bsy_1_1 : 1'b1 ) &&
										( (id == 6'b000100) ? soc1.core.rob.rob_bsy__2 : 1'b1 ) &&
										( (id == 6'b000101) ? soc1.core.rob.rob_bsy_1_2 : 1'b1 ) &&
										( (id == 6'b000110) ? soc1.core.rob.rob_bsy__3 : 1'b1 ) &&
										( (id == 6'b000111) ? soc1.core.rob.rob_bsy_1_3 : 1'b1 ) &&
										( (id == 6'b001000) ? soc1.core.rob.rob_bsy__4 : 1'b1 ) &&
										( (id == 6'b001001) ? soc1.core.rob.rob_bsy_1_4 : 1'b1 ) &&
										( (id == 6'b001010) ? soc1.core.rob.rob_bsy__5 : 1'b1 ) &&
										( (id == 6'b001011) ? soc1.core.rob.rob_bsy_1_5 : 1'b1 ) &&
										( (id == 6'b001100) ? soc1.core.rob.rob_bsy__6 : 1'b1 ) &&
										( (id == 6'b001101) ? soc1.core.rob.rob_bsy_1_6 : 1'b1 ) &&
										( (id == 6'b001110) ? soc1.core.rob.rob_bsy__7 : 1'b1 ) &&
										( (id == 6'b001111) ? soc1.core.rob.rob_bsy_1_7 : 1'b1 ) &&
										( (id == 6'b010000) ? soc1.core.rob.rob_bsy__8 : 1'b1 ) &&
										( (id == 6'b010001) ? soc1.core.rob.rob_bsy_1_8 : 1'b1 ) &&
										( (id == 6'b010010) ? soc1.core.rob.rob_bsy__9 : 1'b1 ) &&
										( (id == 6'b010011) ? soc1.core.rob.rob_bsy_1_9 : 1'b1 ) &&
										( (id == 6'b010100) ? soc1.core.rob.rob_bsy__10 : 1'b1 ) &&
										( (id == 6'b010101) ? soc1.core.rob.rob_bsy_1_10 : 1'b1 ) &&
										( (id == 6'b010110) ? soc1.core.rob.rob_bsy__11 : 1'b1 ) &&
										( (id == 6'b010111) ? soc1.core.rob.rob_bsy_1_11 : 1'b1 ) &&
										( (id == 6'b011000) ? soc1.core.rob.rob_bsy__12 : 1'b1 ) &&
										( (id == 6'b011001) ? soc1.core.rob.rob_bsy_1_12 : 1'b1 ) &&
										( (id == 6'b011010) ? soc1.core.rob.rob_bsy__13 : 1'b1 ) &&
										( (id == 6'b011011) ? soc1.core.rob.rob_bsy_1_13 : 1'b1 ) &&
										( (id == 6'b011100) ? soc1.core.rob.rob_bsy__14 : 1'b1 ) &&
										( (id == 6'b011101) ? soc1.core.rob.rob_bsy_1_14 : 1'b1 ) &&
										( (id == 6'b011110) ? soc1.core.rob.rob_bsy__15 : 1'b1 ) &&
										( (id == 6'b011111) ? soc1.core.rob.rob_bsy_1_15 : 1'b1 ) &&
										( (id == 6'b100000) ? soc1.core.rob.rob_bsy__16 : 1'b1 ) &&
										( (id == 6'b100001) ? soc1.core.rob.rob_bsy_1_16 : 1'b1 ) &&
										( (id == 6'b100010) ? soc1.core.rob.rob_bsy__17 : 1'b1 ) &&
										( (id == 6'b100011) ? soc1.core.rob.rob_bsy_1_17 : 1'b1 ) &&
										( (id == 6'b100100) ? soc1.core.rob.rob_bsy__18 : 1'b1 ) &&
										( (id == 6'b100101) ? soc1.core.rob.rob_bsy_1_18 : 1'b1 ) &&
										( (id == 6'b100110) ? soc1.core.rob.rob_bsy__19 : 1'b1 ) &&
										( (id == 6'b100111) ? soc1.core.rob.rob_bsy_1_19 : 1'b1 ) &&
										( (id == 6'b101000) ? soc1.core.rob.rob_bsy__20 : 1'b1 ) &&
										( (id == 6'b101001) ? soc1.core.rob.rob_bsy_1_20 : 1'b1 ) &&
										( (id == 6'b101010) ? soc1.core.rob.rob_bsy__21 : 1'b1 ) &&
										( (id == 6'b101011) ? soc1.core.rob.rob_bsy_1_21 : 1'b1 ) &&
										( (id == 6'b101100) ? soc1.core.rob.rob_bsy__22 : 1'b1 ) &&
										( (id == 6'b101101) ? soc1.core.rob.rob_bsy_1_22 : 1'b1 ) &&
										( (id == 6'b101110) ? soc1.core.rob.rob_bsy__23 : 1'b1 ) &&
										( (id == 6'b101111) ? soc1.core.rob.rob_bsy_1_23 : 1'b1 ) &&
										( (id == 6'b110000) ? soc1.core.rob.rob_bsy__24 : 1'b1 ) &&
										( (id == 6'b110001) ? soc1.core.rob.rob_bsy_1_24 : 1'b1 ) &&
										( (id == 6'b110010) ? soc1.core.rob.rob_bsy__25 : 1'b1 ) &&
										( (id == 6'b110011) ? soc1.core.rob.rob_bsy_1_25 : 1'b1 ) &&
										( (id == 6'b110100) ? soc1.core.rob.rob_bsy__26 : 1'b1 ) &&
										( (id == 6'b110101) ? soc1.core.rob.rob_bsy_1_26 : 1'b1 ) &&
										( (id == 6'b110110) ? soc1.core.rob.rob_bsy__27 : 1'b1 ) &&
										( (id == 6'b110111) ? soc1.core.rob.rob_bsy_1_27 : 1'b1 ) &&
										( (id == 6'b111000) ? soc1.core.rob.rob_bsy__28 : 1'b1 ) &&
										( (id == 6'b111001) ? soc1.core.rob.rob_bsy_1_28 : 1'b1 ) &&
										( (id == 6'b111010) ? soc1.core.rob.rob_bsy__29 : 1'b1 ) &&
										( (id == 6'b111011) ? soc1.core.rob.rob_bsy_1_29 : 1'b1 ) &&
										( (id == 6'b111100) ? soc1.core.rob.rob_bsy__30 : 1'b1 ) &&
										( (id == 6'b111101) ? soc1.core.rob.rob_bsy_1_30 : 1'b1 ) &&
										( (id == 6'b111110) ? soc1.core.rob.rob_bsy__31 : 1'b1 ) &&
										( (id == 6'b111111) ? soc1.core.rob.rob_bsy_1_31 : 1'b1 );
		end
	endfunction

  //Function that returns if the given ID in the ROB in SoC2 has its busy bit set
	function automatic isPending_2;
		input [5:0] id;
		begin
			isPending_2 = ( (id == 6'b000000) ? soc2.core.rob.rob_bsy__0 : 1'b1 ) &&
										( (id == 6'b000001) ? soc2.core.rob.rob_bsy_1_0 : 1'b1 ) &&
										( (id == 6'b000010) ? soc2.core.rob.rob_bsy__1 : 1'b1 ) &&
										( (id == 6'b000011) ? soc2.core.rob.rob_bsy_1_1 : 1'b1 ) &&
										( (id == 6'b000100) ? soc2.core.rob.rob_bsy__2 : 1'b1 ) &&
										( (id == 6'b000101) ? soc2.core.rob.rob_bsy_1_2 : 1'b1 ) &&
										( (id == 6'b000110) ? soc2.core.rob.rob_bsy__3 : 1'b1 ) &&
										( (id == 6'b000111) ? soc2.core.rob.rob_bsy_1_3 : 1'b1 ) &&
										( (id == 6'b001000) ? soc2.core.rob.rob_bsy__4 : 1'b1 ) &&
										( (id == 6'b001001) ? soc2.core.rob.rob_bsy_1_4 : 1'b1 ) &&
										( (id == 6'b001010) ? soc2.core.rob.rob_bsy__5 : 1'b1 ) &&
										( (id == 6'b001011) ? soc2.core.rob.rob_bsy_1_5 : 1'b1 ) &&
										( (id == 6'b001100) ? soc2.core.rob.rob_bsy__6 : 1'b1 ) &&
										( (id == 6'b001101) ? soc2.core.rob.rob_bsy_1_6 : 1'b1 ) &&
										( (id == 6'b001110) ? soc2.core.rob.rob_bsy__7 : 1'b1 ) &&
										( (id == 6'b001111) ? soc2.core.rob.rob_bsy_1_7 : 1'b1 ) &&
										( (id == 6'b010000) ? soc2.core.rob.rob_bsy__8 : 1'b1 ) &&
										( (id == 6'b010001) ? soc2.core.rob.rob_bsy_1_8 : 1'b1 ) &&
										( (id == 6'b010010) ? soc2.core.rob.rob_bsy__9 : 1'b1 ) &&
										( (id == 6'b010011) ? soc2.core.rob.rob_bsy_1_9 : 1'b1 ) &&
										( (id == 6'b010100) ? soc2.core.rob.rob_bsy__10 : 1'b1 ) &&
										( (id == 6'b010101) ? soc2.core.rob.rob_bsy_1_10 : 1'b1 ) &&
										( (id == 6'b010110) ? soc2.core.rob.rob_bsy__11 : 1'b1 ) &&
										( (id == 6'b010111) ? soc2.core.rob.rob_bsy_1_11 : 1'b1 ) &&
										( (id == 6'b011000) ? soc2.core.rob.rob_bsy__12 : 1'b1 ) &&
										( (id == 6'b011001) ? soc2.core.rob.rob_bsy_1_12 : 1'b1 ) &&
										( (id == 6'b011010) ? soc2.core.rob.rob_bsy__13 : 1'b1 ) &&
										( (id == 6'b011011) ? soc2.core.rob.rob_bsy_1_13 : 1'b1 ) &&
										( (id == 6'b011100) ? soc2.core.rob.rob_bsy__14 : 1'b1 ) &&
										( (id == 6'b011101) ? soc2.core.rob.rob_bsy_1_14 : 1'b1 ) &&
										( (id == 6'b011110) ? soc2.core.rob.rob_bsy__15 : 1'b1 ) &&
										( (id == 6'b011111) ? soc2.core.rob.rob_bsy_1_15 : 1'b1 ) &&
										( (id == 6'b100000) ? soc2.core.rob.rob_bsy__16 : 1'b1 ) &&
										( (id == 6'b100001) ? soc2.core.rob.rob_bsy_1_16 : 1'b1 ) &&
										( (id == 6'b100010) ? soc2.core.rob.rob_bsy__17 : 1'b1 ) &&
										( (id == 6'b100011) ? soc2.core.rob.rob_bsy_1_17 : 1'b1 ) &&
										( (id == 6'b100100) ? soc2.core.rob.rob_bsy__18 : 1'b1 ) &&
										( (id == 6'b100101) ? soc2.core.rob.rob_bsy_1_18 : 1'b1 ) &&
										( (id == 6'b100110) ? soc2.core.rob.rob_bsy__19 : 1'b1 ) &&
										( (id == 6'b100111) ? soc2.core.rob.rob_bsy_1_19 : 1'b1 ) &&
										( (id == 6'b101000) ? soc2.core.rob.rob_bsy__20 : 1'b1 ) &&
										( (id == 6'b101001) ? soc2.core.rob.rob_bsy_1_20 : 1'b1 ) &&
										( (id == 6'b101010) ? soc2.core.rob.rob_bsy__21 : 1'b1 ) &&
										( (id == 6'b101011) ? soc2.core.rob.rob_bsy_1_21 : 1'b1 ) &&
										( (id == 6'b101100) ? soc2.core.rob.rob_bsy__22 : 1'b1 ) &&
										( (id == 6'b101101) ? soc2.core.rob.rob_bsy_1_22 : 1'b1 ) &&
										( (id == 6'b101110) ? soc2.core.rob.rob_bsy__23 : 1'b1 ) &&
										( (id == 6'b101111) ? soc2.core.rob.rob_bsy_1_23 : 1'b1 ) &&
										( (id == 6'b110000) ? soc2.core.rob.rob_bsy__24 : 1'b1 ) &&
										( (id == 6'b110001) ? soc2.core.rob.rob_bsy_1_24 : 1'b1 ) &&
										( (id == 6'b110010) ? soc2.core.rob.rob_bsy__25 : 1'b1 ) &&
										( (id == 6'b110011) ? soc2.core.rob.rob_bsy_1_25 : 1'b1 ) &&
										( (id == 6'b110100) ? soc2.core.rob.rob_bsy__26 : 1'b1 ) &&
										( (id == 6'b110101) ? soc2.core.rob.rob_bsy_1_26 : 1'b1 ) &&
										( (id == 6'b110110) ? soc2.core.rob.rob_bsy__27 : 1'b1 ) &&
										( (id == 6'b110111) ? soc2.core.rob.rob_bsy_1_27 : 1'b1 ) &&
										( (id == 6'b111000) ? soc2.core.rob.rob_bsy__28 : 1'b1 ) &&
										( (id == 6'b111001) ? soc2.core.rob.rob_bsy_1_28 : 1'b1 ) &&
										( (id == 6'b111010) ? soc2.core.rob.rob_bsy__29 : 1'b1 ) &&
										( (id == 6'b111011) ? soc2.core.rob.rob_bsy_1_29 : 1'b1 ) &&
										( (id == 6'b111100) ? soc2.core.rob.rob_bsy__30 : 1'b1 ) &&
										( (id == 6'b111101) ? soc2.core.rob.rob_bsy_1_30 : 1'b1 ) &&
										( (id == 6'b111110) ? soc2.core.rob.rob_bsy__31 : 1'b1 ) &&
										( (id == 6'b111111) ? soc2.core.rob.rob_bsy_1_31 : 1'b1 );
		end
	endfunction

  //Function that returns if the given ID in the ROB in SoC1 has its valid bit set
	function automatic isValid_1;
		input [5:0] id;
		begin
			isValid_1 = ( (id == 6'b000000) ? soc1.core.rob.rob_val__0 : 1'b1 ) &&
										( (id == 6'b000001) ? soc1.core.rob.rob_val_1_0 : 1'b1 ) &&
										( (id == 6'b000010) ? soc1.core.rob.rob_val__1 : 1'b1 ) &&
										( (id == 6'b000011) ? soc1.core.rob.rob_val_1_1 : 1'b1 ) &&
										( (id == 6'b000100) ? soc1.core.rob.rob_val__2 : 1'b1 ) &&
										( (id == 6'b000101) ? soc1.core.rob.rob_val_1_2 : 1'b1 ) &&
										( (id == 6'b000110) ? soc1.core.rob.rob_val__3 : 1'b1 ) &&
										( (id == 6'b000111) ? soc1.core.rob.rob_val_1_3 : 1'b1 ) &&
										( (id == 6'b001000) ? soc1.core.rob.rob_val__4 : 1'b1 ) &&
										( (id == 6'b001001) ? soc1.core.rob.rob_val_1_4 : 1'b1 ) &&
										( (id == 6'b001010) ? soc1.core.rob.rob_val__5 : 1'b1 ) &&
										( (id == 6'b001011) ? soc1.core.rob.rob_val_1_5 : 1'b1 ) &&
										( (id == 6'b001100) ? soc1.core.rob.rob_val__6 : 1'b1 ) &&
										( (id == 6'b001101) ? soc1.core.rob.rob_val_1_6 : 1'b1 ) &&
										( (id == 6'b001110) ? soc1.core.rob.rob_val__7 : 1'b1 ) &&
										( (id == 6'b001111) ? soc1.core.rob.rob_val_1_7 : 1'b1 ) &&
										( (id == 6'b010000) ? soc1.core.rob.rob_val__8 : 1'b1 ) &&
										( (id == 6'b010001) ? soc1.core.rob.rob_val_1_8 : 1'b1 ) &&
										( (id == 6'b010010) ? soc1.core.rob.rob_val__9 : 1'b1 ) &&
										( (id == 6'b010011) ? soc1.core.rob.rob_val_1_9 : 1'b1 ) &&
										( (id == 6'b010100) ? soc1.core.rob.rob_val__10 : 1'b1 ) &&
										( (id == 6'b010101) ? soc1.core.rob.rob_val_1_10 : 1'b1 ) &&
										( (id == 6'b010110) ? soc1.core.rob.rob_val__11 : 1'b1 ) &&
										( (id == 6'b010111) ? soc1.core.rob.rob_val_1_11 : 1'b1 ) &&
										( (id == 6'b011000) ? soc1.core.rob.rob_val__12 : 1'b1 ) &&
										( (id == 6'b011001) ? soc1.core.rob.rob_val_1_12 : 1'b1 ) &&
										( (id == 6'b011010) ? soc1.core.rob.rob_val__13 : 1'b1 ) &&
										( (id == 6'b011011) ? soc1.core.rob.rob_val_1_13 : 1'b1 ) &&
										( (id == 6'b011100) ? soc1.core.rob.rob_val__14 : 1'b1 ) &&
										( (id == 6'b011101) ? soc1.core.rob.rob_val_1_14 : 1'b1 ) &&
										( (id == 6'b011110) ? soc1.core.rob.rob_val__15 : 1'b1 ) &&
										( (id == 6'b011111) ? soc1.core.rob.rob_val_1_15 : 1'b1 ) &&
										( (id == 6'b100000) ? soc1.core.rob.rob_val__16 : 1'b1 ) &&
										( (id == 6'b100001) ? soc1.core.rob.rob_val_1_16 : 1'b1 ) &&
										( (id == 6'b100010) ? soc1.core.rob.rob_val__17 : 1'b1 ) &&
										( (id == 6'b100011) ? soc1.core.rob.rob_val_1_17 : 1'b1 ) &&
										( (id == 6'b100100) ? soc1.core.rob.rob_val__18 : 1'b1 ) &&
										( (id == 6'b100101) ? soc1.core.rob.rob_val_1_18 : 1'b1 ) &&
										( (id == 6'b100110) ? soc1.core.rob.rob_val__19 : 1'b1 ) &&
										( (id == 6'b100111) ? soc1.core.rob.rob_val_1_19 : 1'b1 ) &&
										( (id == 6'b101000) ? soc1.core.rob.rob_val__20 : 1'b1 ) &&
										( (id == 6'b101001) ? soc1.core.rob.rob_val_1_20 : 1'b1 ) &&
										( (id == 6'b101010) ? soc1.core.rob.rob_val__21 : 1'b1 ) &&
										( (id == 6'b101011) ? soc1.core.rob.rob_val_1_21 : 1'b1 ) &&
										( (id == 6'b101100) ? soc1.core.rob.rob_val__22 : 1'b1 ) &&
										( (id == 6'b101101) ? soc1.core.rob.rob_val_1_22 : 1'b1 ) &&
										( (id == 6'b101110) ? soc1.core.rob.rob_val__23 : 1'b1 ) &&
										( (id == 6'b101111) ? soc1.core.rob.rob_val_1_23 : 1'b1 ) &&
										( (id == 6'b110000) ? soc1.core.rob.rob_val__24 : 1'b1 ) &&
										( (id == 6'b110001) ? soc1.core.rob.rob_val_1_24 : 1'b1 ) &&
										( (id == 6'b110010) ? soc1.core.rob.rob_val__25 : 1'b1 ) &&
										( (id == 6'b110011) ? soc1.core.rob.rob_val_1_25 : 1'b1 ) &&
										( (id == 6'b110100) ? soc1.core.rob.rob_val__26 : 1'b1 ) &&
										( (id == 6'b110101) ? soc1.core.rob.rob_val_1_26 : 1'b1 ) &&
										( (id == 6'b110110) ? soc1.core.rob.rob_val__27 : 1'b1 ) &&
										( (id == 6'b110111) ? soc1.core.rob.rob_val_1_27 : 1'b1 ) &&
										( (id == 6'b111000) ? soc1.core.rob.rob_val__28 : 1'b1 ) &&
										( (id == 6'b111001) ? soc1.core.rob.rob_val_1_28 : 1'b1 ) &&
										( (id == 6'b111010) ? soc1.core.rob.rob_val__29 : 1'b1 ) &&
										( (id == 6'b111011) ? soc1.core.rob.rob_val_1_29 : 1'b1 ) &&
										( (id == 6'b111100) ? soc1.core.rob.rob_val__30 : 1'b1 ) &&
										( (id == 6'b111101) ? soc1.core.rob.rob_val_1_30 : 1'b1 ) &&
										( (id == 6'b111110) ? soc1.core.rob.rob_val__31 : 1'b1 ) &&
										( (id == 6'b111111) ? soc1.core.rob.rob_val_1_31 : 1'b1 );
		end
	endfunction

  //Function that returns if the given ID in the ROB in SoC2 has its busy bit set
	function automatic isValid_2;
		input [5:0] id;
		begin
			isValid_2 = ( (id == 6'b000000) ? soc2.core.rob.rob_val__0 : 1'b1 ) &&
										( (id == 6'b000001) ? soc2.core.rob.rob_val_1_0 : 1'b1 ) &&
										( (id == 6'b000010) ? soc2.core.rob.rob_val__1 : 1'b1 ) &&
										( (id == 6'b000011) ? soc2.core.rob.rob_val_1_1 : 1'b1 ) &&
										( (id == 6'b000100) ? soc2.core.rob.rob_val__2 : 1'b1 ) &&
										( (id == 6'b000101) ? soc2.core.rob.rob_val_1_2 : 1'b1 ) &&
										( (id == 6'b000110) ? soc2.core.rob.rob_val__3 : 1'b1 ) &&
										( (id == 6'b000111) ? soc2.core.rob.rob_val_1_3 : 1'b1 ) &&
										( (id == 6'b001000) ? soc2.core.rob.rob_val__4 : 1'b1 ) &&
										( (id == 6'b001001) ? soc2.core.rob.rob_val_1_4 : 1'b1 ) &&
										( (id == 6'b001010) ? soc2.core.rob.rob_val__5 : 1'b1 ) &&
										( (id == 6'b001011) ? soc2.core.rob.rob_val_1_5 : 1'b1 ) &&
										( (id == 6'b001100) ? soc2.core.rob.rob_val__6 : 1'b1 ) &&
										( (id == 6'b001101) ? soc2.core.rob.rob_val_1_6 : 1'b1 ) &&
										( (id == 6'b001110) ? soc2.core.rob.rob_val__7 : 1'b1 ) &&
										( (id == 6'b001111) ? soc2.core.rob.rob_val_1_7 : 1'b1 ) &&
										( (id == 6'b010000) ? soc2.core.rob.rob_val__8 : 1'b1 ) &&
										( (id == 6'b010001) ? soc2.core.rob.rob_val_1_8 : 1'b1 ) &&
										( (id == 6'b010010) ? soc2.core.rob.rob_val__9 : 1'b1 ) &&
										( (id == 6'b010011) ? soc2.core.rob.rob_val_1_9 : 1'b1 ) &&
										( (id == 6'b010100) ? soc2.core.rob.rob_val__10 : 1'b1 ) &&
										( (id == 6'b010101) ? soc2.core.rob.rob_val_1_10 : 1'b1 ) &&
										( (id == 6'b010110) ? soc2.core.rob.rob_val__11 : 1'b1 ) &&
										( (id == 6'b010111) ? soc2.core.rob.rob_val_1_11 : 1'b1 ) &&
										( (id == 6'b011000) ? soc2.core.rob.rob_val__12 : 1'b1 ) &&
										( (id == 6'b011001) ? soc2.core.rob.rob_val_1_12 : 1'b1 ) &&
										( (id == 6'b011010) ? soc2.core.rob.rob_val__13 : 1'b1 ) &&
										( (id == 6'b011011) ? soc2.core.rob.rob_val_1_13 : 1'b1 ) &&
										( (id == 6'b011100) ? soc2.core.rob.rob_val__14 : 1'b1 ) &&
										( (id == 6'b011101) ? soc2.core.rob.rob_val_1_14 : 1'b1 ) &&
										( (id == 6'b011110) ? soc2.core.rob.rob_val__15 : 1'b1 ) &&
										( (id == 6'b011111) ? soc2.core.rob.rob_val_1_15 : 1'b1 ) &&
										( (id == 6'b100000) ? soc2.core.rob.rob_val__16 : 1'b1 ) &&
										( (id == 6'b100001) ? soc2.core.rob.rob_val_1_16 : 1'b1 ) &&
										( (id == 6'b100010) ? soc2.core.rob.rob_val__17 : 1'b1 ) &&
										( (id == 6'b100011) ? soc2.core.rob.rob_val_1_17 : 1'b1 ) &&
										( (id == 6'b100100) ? soc2.core.rob.rob_val__18 : 1'b1 ) &&
										( (id == 6'b100101) ? soc2.core.rob.rob_val_1_18 : 1'b1 ) &&
										( (id == 6'b100110) ? soc2.core.rob.rob_val__19 : 1'b1 ) &&
										( (id == 6'b100111) ? soc2.core.rob.rob_val_1_19 : 1'b1 ) &&
										( (id == 6'b101000) ? soc2.core.rob.rob_val__20 : 1'b1 ) &&
										( (id == 6'b101001) ? soc2.core.rob.rob_val_1_20 : 1'b1 ) &&
										( (id == 6'b101010) ? soc2.core.rob.rob_val__21 : 1'b1 ) &&
										( (id == 6'b101011) ? soc2.core.rob.rob_val_1_21 : 1'b1 ) &&
										( (id == 6'b101100) ? soc2.core.rob.rob_val__22 : 1'b1 ) &&
										( (id == 6'b101101) ? soc2.core.rob.rob_val_1_22 : 1'b1 ) &&
										( (id == 6'b101110) ? soc2.core.rob.rob_val__23 : 1'b1 ) &&
										( (id == 6'b101111) ? soc2.core.rob.rob_val_1_23 : 1'b1 ) &&
										( (id == 6'b110000) ? soc2.core.rob.rob_val__24 : 1'b1 ) &&
										( (id == 6'b110001) ? soc2.core.rob.rob_val_1_24 : 1'b1 ) &&
										( (id == 6'b110010) ? soc2.core.rob.rob_val__25 : 1'b1 ) &&
										( (id == 6'b110011) ? soc2.core.rob.rob_val_1_25 : 1'b1 ) &&
										( (id == 6'b110100) ? soc2.core.rob.rob_val__26 : 1'b1 ) &&
										( (id == 6'b110101) ? soc2.core.rob.rob_val_1_26 : 1'b1 ) &&
										( (id == 6'b110110) ? soc2.core.rob.rob_val__27 : 1'b1 ) &&
										( (id == 6'b110111) ? soc2.core.rob.rob_val_1_27 : 1'b1 ) &&
										( (id == 6'b111000) ? soc2.core.rob.rob_val__28 : 1'b1 ) &&
										( (id == 6'b111001) ? soc2.core.rob.rob_val_1_28 : 1'b1 ) &&
										( (id == 6'b111010) ? soc2.core.rob.rob_val__29 : 1'b1 ) &&
										( (id == 6'b111011) ? soc2.core.rob.rob_val_1_29 : 1'b1 ) &&
										( (id == 6'b111100) ? soc2.core.rob.rob_val__30 : 1'b1 ) &&
										( (id == 6'b111101) ? soc2.core.rob.rob_val_1_30 : 1'b1 ) &&
										( (id == 6'b111110) ? soc2.core.rob.rob_val__31 : 1'b1 ) &&
										( (id == 6'b111111) ? soc2.core.rob.rob_val_1_31 : 1'b1 );
		end
	endfunction

  //Function that returns if the given row is in the committable set
  //to be committable, the ID of the row must be above head and below or equal to root_id
	function automatic isRobRowCommitable;
		input [4:0] head_id;
		input [5:0] root_id;
		input [4:0] row;
		begin
      //since the ROB is a ringbuffer, we need to distinguish different cases for the position of head and root_id
			if (head_id < root_id[5:1])
			begin
				isRobRowCommitable =  row >= head_id && row < root_id[5:1];
			end
			else if (head_id > root_id[5:1])
			begin
				isRobRowCommitable = row >= head_id || row < root_id[5:1];
			end
			else // head_id == root_id
			begin
				isRobRowCommitable = ( row == head_id ); // there is no commitable, except for head_id
			end
		end
	endfunction

  //Function that returns if the given ID is in the committable set
  //to be committable, the ID must be above head and below or equal to root_id
	function automatic isRobIdCommitable;
		input [4:0] head_id;
		input [5:0] root_id;
		input [5:0] id;
		begin
      //since the ROB is a ringbuffer, we need to distinguish different cases for the position of head and root_id
			if (head_id < root_id[5:1])
			begin
				isRobIdCommitable =  id[5:1] >= head_id && id <= root_id;
			end
			else if (head_id > root_id[5:1])
			begin
				isRobIdCommitable = id[5:1] >= head_id || id <= root_id;
			end
			else // head_id == root_id
			begin
				isRobIdCommitable = ( id == root_id ); // there is no commitable, except for root_id
			end

		end
	endfunction

  //function that returns true if the given spawn_tag is greater than T_main
	function automatic isSpawnTagGreater;
    //4-bit branch tag(spawn_tag), which is the integer value of the level of speculation
		input [3:0] spawn_tag;
		input [11:0] main_tag;
		reg [15:0] temp;
		reg [11:0] temp2;
		begin
      //constructs a 12-bit branch mask by shifting a 1 by the value of the branch tag
			temp = (16'h1 << spawn_tag);
			temp2 = temp[11:0];
      //check if the intersection of the branch mask and the main_tag (T_main) is 0
      //then the spawn_tag is greater than T_main
			isSpawnTagGreater = (temp2 & main_tag) == 12'h0;
		end
	endfunction

//*******************************************//

	wire [5:0] root_id;
	assign root_id = 6'b010000; // should be symbolic

	wire [11:0] root_br_mask; // should be symbolic // let's assume it is onehot
	assign root_br_mask = 12'h080;

  //needed signals for misprediction of instruction at root_id
  //see template for more information
	reg mispred_flag_1;
	reg mispred_happened_1;
	reg mispred_flag_2;
	reg mispred_happened_2;

  //combinational logic for setting the flags
	always @(posedge clock)
	begin
		if (reset)
		begin
			mispred_flag_1 <= 1'b0;
			mispred_happened_1 <= 1'b0;
			mispred_flag_2 <= 1'b0;
			mispred_happened_2 <= 1'b0;
		end
		else
		begin
		      //if masks match set the flags
		      if (((soc1.core.rob.io_brupdate_b1_mispredict_mask & rob_branch_masks_1[root_id]) != 12'h0 ||
		      !((soc1.core.rob.rob_head < soc1.core.rob.rob_tail) && (soc1.core.rob.rob_head <= root_id[5:1]) && (root_id[5:1] < soc1.core.rob.rob_tail)
		      ||
		      !(soc1.core.rob.rob_head < soc1.core.rob.rob_tail) && (soc1.core.rob.rob_head > soc1.core.rob.rob_tail) && ((soc1.core.rob.rob_head <= root_id[5:1]) || (root_id[5:1] < soc1.core.rob.rob_tail))
		      ||
		      !(soc1.core.rob.rob_head < soc1.core.rob.rob_tail) && !(soc1.core.rob.rob_head > soc1.core.rob.rob_tail) && !soc1.core.rob.io_empty )) &&
		     	mispred_happened_1 == 1'b0 )
			begin
				mispred_flag_1 <= 1'b1;
				mispred_happened_1 <= 1'b1;
			end
			else
			begin
        			//unset this flag after one clock cycle
				mispred_flag_1 <= 1'b0;
			end

		      //if masks match set the flags
		      if (((soc2.core.rob.io_brupdate_b1_mispredict_mask & rob_branch_masks_2[root_id]) != 12'h0 ||
		      !((soc2.core.rob.rob_head < soc2.core.rob.rob_tail) && (soc2.core.rob.rob_head <= root_id[5:1]) && (root_id[5:1] < soc2.core.rob.rob_tail)
		      ||
		      !(soc2.core.rob.rob_head < soc2.core.rob.rob_tail) && (soc2.core.rob.rob_head > soc2.core.rob.rob_tail) && ((soc2.core.rob.rob_head <= root_id[5:1]) || (root_id[5:1] < soc2.core.rob.rob_tail))
		      ||
		      !(soc2.core.rob.rob_head < soc2.core.rob.rob_tail) && !(soc2.core.rob.rob_head > soc2.core.rob.rob_tail) && !soc2.core.rob.io_empty )) &&
		     	mispred_happened_2 == 1'b0 )
		      begin
				mispred_flag_2 <= 1'b1;
				mispred_happened_2 <= 1'b1;
			end
			else
			begin
        			//unset this flag after one clock cycle
				mispred_flag_2 <= 1'b0;
			end

		end
	end

//****************************************************//
//************ME-1(Main Branch Pending)***************//

  //i) ROB slot with root_ID contains an SPI Instruction
	wire ME_1_1;
  //call to isSpi function
	assign ME_1_1 = (mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed) ? isSpi(root_id) : 1'b1;

  //ii) SPI is mispredicted
	wire ME_1_2;
  //SPI is mispredicted if it is never correct predicted
	assign ME_1_2 = ( (mispred_happened_1 == 1'b0) && (!root_id_killed && !root_id_already_killed) && soc1.core.brinfos_0_valid && !soc1.core.brinfos_0_mispredict ? soc1.core.brinfos_0_uop_br_tag != 4'h7 : 1'b1 ) &&
                  ( (mispred_happened_1 == 1'b0) && (!root_id_killed && !root_id_already_killed) && soc1.core.brinfos_1_valid && !soc1.core.brinfos_1_mispredict ? soc1.core.brinfos_1_uop_br_tag != 4'h7 : 1'b1 ) &&
                  ( (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed) && soc2.core.brinfos_0_valid && !soc2.core.brinfos_0_mispredict ? soc2.core.brinfos_0_uop_br_tag != 4'h7 : 1'b1 ) &&
                  ( (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed) && soc2.core.brinfos_1_valid && !soc2.core.brinfos_1_mispredict ? soc2.core.brinfos_1_uop_br_tag != 4'h7 : 1'b1 );

  //iii) SPI remains valid(pending) until misprediction is signaled by the prediction unit
	wire ME_1_3;
  // check busy and valid bit
  assign ME_1_3 = ( (mispred_happened_1 == 1'b0) && (!root_id_killed && !root_id_already_killed) ? isPending_1(root_id) && isValid_1(root_id) : 1'b1 ) && ( (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed) ? isPending_2(root_id) && isValid_2(root_id) : 1'b1 );

	wire ME_1;
	assign ME_1 = ME_1_1 && ME_1_2 && ME_1_3;


//****************************************************//
//************ME-2(Uncommittable Slots Invalidated)***//

	wire ME_2_1;
  //after misprediction of SPI, in the next clock cycle every ROB slot in the uncommittable set is invalidated (SoC1)
	assign ME_2_1 = (mispred_flag_1 && (soc1.core.rob.rob_state != 2'h2)) && (!root_id_killed && !root_id_already_killed) ? ( ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000000 ) || soc1.core.rob.rob_val__0 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000001 ) || soc1.core.rob.rob_val_1_0 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000010 ) || soc1.core.rob.rob_val__1 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000011 ) || soc1.core.rob.rob_val_1_1 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000100 ) || soc1.core.rob.rob_val__2 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000101 ) || soc1.core.rob.rob_val_1_2 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000110 ) || soc1.core.rob.rob_val__3 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000111 ) || soc1.core.rob.rob_val_1_3 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001000 ) || soc1.core.rob.rob_val__4 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001001 ) || soc1.core.rob.rob_val_1_4 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001010 ) || soc1.core.rob.rob_val__5 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001011 ) || soc1.core.rob.rob_val_1_5 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001100 ) || soc1.core.rob.rob_val__6 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001101 ) || soc1.core.rob.rob_val_1_6 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001110 ) || soc1.core.rob.rob_val__7 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001111 ) || soc1.core.rob.rob_val_1_7 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010000 ) || soc1.core.rob.rob_val__8 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010001 ) || soc1.core.rob.rob_val_1_8 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010010 ) || soc1.core.rob.rob_val__9 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010011 ) || soc1.core.rob.rob_val_1_9 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010100 ) || soc1.core.rob.rob_val__10 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010101 ) || soc1.core.rob.rob_val_1_10 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010110 ) || soc1.core.rob.rob_val__11 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010111 ) || soc1.core.rob.rob_val_1_11 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011000 ) || soc1.core.rob.rob_val__12 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011001 ) || soc1.core.rob.rob_val_1_12 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011010 ) || soc1.core.rob.rob_val__13 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011011 ) || soc1.core.rob.rob_val_1_13 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011100 ) || soc1.core.rob.rob_val__14 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011101 ) || soc1.core.rob.rob_val_1_14 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011110 ) || soc1.core.rob.rob_val__15 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011111 ) || soc1.core.rob.rob_val_1_15 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100000 ) || soc1.core.rob.rob_val__16 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100001 ) || soc1.core.rob.rob_val_1_16 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100010 ) || soc1.core.rob.rob_val__17 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100011 ) || soc1.core.rob.rob_val_1_17 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100100 ) || soc1.core.rob.rob_val__18 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100101 ) || soc1.core.rob.rob_val_1_18 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100110 ) || soc1.core.rob.rob_val__19 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100111 ) || soc1.core.rob.rob_val_1_19 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101000 ) || soc1.core.rob.rob_val__20 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101001 ) || soc1.core.rob.rob_val_1_20 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101010 ) || soc1.core.rob.rob_val__21 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101011 ) || soc1.core.rob.rob_val_1_21 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101100 ) || soc1.core.rob.rob_val__22 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101101 ) || soc1.core.rob.rob_val_1_22 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101110 ) || soc1.core.rob.rob_val__23 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101111 ) || soc1.core.rob.rob_val_1_23 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110000 ) || soc1.core.rob.rob_val__24 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110001 ) || soc1.core.rob.rob_val_1_24 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110010 ) || soc1.core.rob.rob_val__25 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110011 ) || soc1.core.rob.rob_val_1_25 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110100 ) || soc1.core.rob.rob_val__26 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110101 ) || soc1.core.rob.rob_val_1_26 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110110 ) || soc1.core.rob.rob_val__27 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110111 ) || soc1.core.rob.rob_val_1_27 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111000 ) || soc1.core.rob.rob_val__28 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111001 ) || soc1.core.rob.rob_val_1_28 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111010 ) || soc1.core.rob.rob_val__29 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111011 ) || soc1.core.rob.rob_val_1_29 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111100 ) || soc1.core.rob.rob_val__30 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111101 ) || soc1.core.rob.rob_val_1_30 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111110 ) || soc1.core.rob.rob_val__31 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111111 ) || soc1.core.rob.rob_val_1_31 == 1'b0 )
																			) : 1'b1;

	wire ME_2_2;
  //after misprediction of SPI, in the next clock cycle every ROB slot in the uncommittable set is invalidated (SoC2)
	assign ME_2_2 = (mispred_flag_2 && (soc2.core.rob.rob_state != 2'h2)) && (!root_id_killed && !root_id_already_killed) ? ( ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000000 ) || soc2.core.rob.rob_val__0 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000001 ) || soc2.core.rob.rob_val_1_0 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000010 ) || soc2.core.rob.rob_val__1 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000011 ) || soc2.core.rob.rob_val_1_1 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000100 ) || soc2.core.rob.rob_val__2 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000101 ) || soc2.core.rob.rob_val_1_2 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000110 ) || soc2.core.rob.rob_val__3 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000111 ) || soc2.core.rob.rob_val_1_3 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001000 ) || soc2.core.rob.rob_val__4 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001001 ) || soc2.core.rob.rob_val_1_4 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001010 ) || soc2.core.rob.rob_val__5 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001011 ) || soc2.core.rob.rob_val_1_5 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001100 ) || soc2.core.rob.rob_val__6 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001101 ) || soc2.core.rob.rob_val_1_6 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001110 ) || soc2.core.rob.rob_val__7 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001111 ) || soc2.core.rob.rob_val_1_7 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010000 ) || soc2.core.rob.rob_val__8 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010001 ) || soc2.core.rob.rob_val_1_8 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010010 ) || soc2.core.rob.rob_val__9 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010011 ) || soc2.core.rob.rob_val_1_9 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010100 ) || soc2.core.rob.rob_val__10 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010101 ) || soc2.core.rob.rob_val_1_10 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010110 ) || soc2.core.rob.rob_val__11 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010111 ) || soc2.core.rob.rob_val_1_11 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011000 ) || soc2.core.rob.rob_val__12 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011001 ) || soc2.core.rob.rob_val_1_12 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011010 ) || soc2.core.rob.rob_val__13 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011011 ) || soc2.core.rob.rob_val_1_13 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011100 ) || soc2.core.rob.rob_val__14 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011101 ) || soc2.core.rob.rob_val_1_14 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011110 ) || soc2.core.rob.rob_val__15 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011111 ) || soc2.core.rob.rob_val_1_15 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100000 ) || soc2.core.rob.rob_val__16 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100001 ) || soc2.core.rob.rob_val_1_16 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100010 ) || soc2.core.rob.rob_val__17 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100011 ) || soc2.core.rob.rob_val_1_17 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100100 ) || soc2.core.rob.rob_val__18 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100101 ) || soc2.core.rob.rob_val_1_18 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100110 ) || soc2.core.rob.rob_val__19 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100111 ) || soc2.core.rob.rob_val_1_19 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101000 ) || soc2.core.rob.rob_val__20 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101001 ) || soc2.core.rob.rob_val_1_20 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101010 ) || soc2.core.rob.rob_val__21 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101011 ) || soc2.core.rob.rob_val_1_21 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101100 ) || soc2.core.rob.rob_val__22 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101101 ) || soc2.core.rob.rob_val_1_22 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101110 ) || soc2.core.rob.rob_val__23 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101111 ) || soc2.core.rob.rob_val_1_23 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110000 ) || soc2.core.rob.rob_val__24 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110001 ) || soc2.core.rob.rob_val_1_24 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110010 ) || soc2.core.rob.rob_val__25 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110011 ) || soc2.core.rob.rob_val_1_25 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110100 ) || soc2.core.rob.rob_val__26 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110101 ) || soc2.core.rob.rob_val_1_26 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110110 ) || soc2.core.rob.rob_val__27 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110111 ) || soc2.core.rob.rob_val_1_27 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111000 ) || soc2.core.rob.rob_val__28 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111001 ) || soc2.core.rob.rob_val_1_28 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111010 ) || soc2.core.rob.rob_val__29 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111011 ) || soc2.core.rob.rob_val_1_29 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111100 ) || soc2.core.rob.rob_val__30 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111101 ) || soc2.core.rob.rob_val_1_30 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111110 ) || soc2.core.rob.rob_val__31 == 1'b0 ) &&
																			 ( isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111111 ) || soc2.core.rob.rob_val_1_31 == 1'b0 )
																			) : 1'b1;

	wire ME_2;
	assign ME_2 = ME_2_1 && ME_2_2;

//****************************************************//
//************ME-3(ROB tail Consistency)**************//

	wire ME_3;
  //until misprediction, ROB tail points to an uncommittable ROB slot
	assign ME_3 = ( (mispred_happened_1 == 1'b0) && (!root_id_killed && !root_id_already_killed) ? ( isRobRowCommitable(soc1.core.rob.rob_head, root_id, soc1.core.rob.rob_tail) == 1'b0 ) : 1'b1 ) &&
								( (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed) ? ( isRobRowCommitable(soc2.core.rob.rob_head, root_id, soc2.core.rob.rob_tail) == 1'b0 ) : 1'b1 )
                ||
                //if head == tail, ROB is either full or empty
                //in both cases, tail does not have to point to an uncommitable slot
                (soc1.core.rob.rob_head == soc1.core.rob.rob_tail) &&
                (soc2.core.rob.rob_head == soc2.core.rob.rob_tail);

//****************************************************//
//************ME-4(FU Consistency))*******************//
//Should we check for request valid bit?
//check for every FU:
//if ROB_IDs of the instructions currently being executed are equal, and commitable,
//the operands must be equal

	wire ME_4_alu;
	assign ME_4_alu = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
                      soc1.core.csr_exe_unit.alu.io_req_bits_uop_rob_idx == soc2.core.csr_exe_unit.alu.io_req_bits_uop_rob_idx &&
										(  soc1.core.csr_exe_unit.alu.io_req_bits_rs1_data != soc2.core.csr_exe_unit.alu.io_req_bits_rs1_data ||
												soc1.core.csr_exe_unit.alu.io_req_bits_rs2_data != soc2.core.csr_exe_unit.alu.io_req_bits_rs2_data ) ) ?
												 isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.csr_exe_unit.alu.io_req_bits_uop_rob_idx) == 1'b0 : 1'b1;

	wire ME_4_div;
	assign ME_4_div = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) && */
                      soc1.core.csr_exe_unit.div.io_req_bits_uop_rob_idx == soc2.core.csr_exe_unit.div.io_req_bits_uop_rob_idx &&
										 ( soc1.core.csr_exe_unit.div.io_req_bits_rs1_data != soc2.core.csr_exe_unit.div.io_req_bits_rs1_data ||
										  soc1.core.csr_exe_unit.div.io_req_bits_rs2_data != soc2.core.csr_exe_unit.div.io_req_bits_rs2_data ) ) ?
											 !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.csr_exe_unit.div.io_req_bits_uop_rob_idx) &&
											 !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.csr_exe_unit.div.io_req_bits_uop_yrot)											 
											 : 1'b1;


  wire ME_4_fpiu;
  assign ME_4_fpiu =  (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
    soc1.core.fp_pipeline.fpiu_unit.io_req_bits_uop_rob_idx == soc2.core.fp_pipeline.fpiu_unit.io_req_bits_uop_rob_idx &&
 ( soc1.core.fp_pipeline.fpiu_unit.io_req_bits_rs1_data != soc2.core.fp_pipeline.fpiu_unit.io_req_bits_rs1_data ||
   soc1.core.fp_pipeline.fpiu_unit.io_req_bits_rs2_data != soc2.core.fp_pipeline.fpiu_unit.io_req_bits_rs2_data ||
   soc1.core.fp_pipeline.fpiu_unit.io_req_bits_rs3_data != soc2.core.fp_pipeline.fpiu_unit.io_req_bits_rs3_data ) ) ?
	 isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.io_req_bits_uop_rob_idx) == 1'b0 : 1'b1;


  wire ME_4_jmpalu;
  assign ME_4_jmpalu =  (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
    soc1.core.jmp_unit.alu.io_req_bits_uop_rob_idx == soc2.core.jmp_unit.alu.io_req_bits_uop_rob_idx &&
 ( soc1.core.jmp_unit.alu.io_req_bits_rs1_data != soc2.core.jmp_unit.alu.io_req_bits_rs1_data ||
   soc1.core.jmp_unit.alu.io_req_bits_rs2_data != soc2.core.jmp_unit.alu.io_req_bits_rs2_data ) ) ?
   !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.alu.io_req_bits_uop_rob_idx) &&
   !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.alu.io_req_bits_uop_yrot)
   : 1'b1;


  wire ME_4_ifpu;
  assign ME_4_ifpu =  (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
    soc1.core.jmp_unit.ifpu.io_req_bits_uop_rob_idx == soc2.core.jmp_unit.ifpu.io_req_bits_uop_rob_idx &&
 ( soc1.core.jmp_unit.ifpu.io_req_bits_rs1_data != soc2.core.jmp_unit.ifpu.io_req_bits_rs1_data ) ) ?
   isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.ifpu.io_req_bits_uop_rob_idx) == 1'b0 : 1'b1;


  wire ME_4_imul;
  assign ME_4_imul =  (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
    soc1.core.jmp_unit.imul.io_req_bits_uop_rob_idx == soc2.core.jmp_unit.imul.io_req_bits_uop_rob_idx &&
 ( soc1.core.jmp_unit.imul.io_req_bits_rs1_data != soc2.core.jmp_unit.imul.io_req_bits_rs1_data ||
   soc1.core.jmp_unit.imul.io_req_bits_rs2_data != soc2.core.jmp_unit.imul.io_req_bits_rs2_data ) ) ?
   isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.imul.io_req_bits_uop_rob_idx) == 1'b0 : 1'b1;


	wire ME_4_lsu;
	assign ME_4_lsu = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
                      soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx == soc2.lsu.io_core_exe_0_req_bits_uop_rob_idx &&
										( soc1.lsu.io_core_exe_0_req_bits_addr != soc2.lsu.io_core_exe_0_req_bits_addr ||
											soc1.lsu.io_core_exe_0_req_bits_data != soc2.lsu.io_core_exe_0_req_bits_data ) )
                      ?
  											(isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx) == 1'b0) &&

                        ((soc1.lsu.io_core_exe_0_req_bits_uop_uses_ldq == 1'b1)
                        ?
                          (
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h0 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_0_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h1 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_1_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h2 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_2_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h3 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_3_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h4 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_4_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h5 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_5_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h6 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_6_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h7 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_7_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h8 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_8_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h9 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_9_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'hb ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_11_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'ha ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_10_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'hc ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_12_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'hd ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_13_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'he ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_14_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'hf ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_15_bits_uop_rob_idx) : 1'b1)
                          )
                        :
                        1'b1)&&

                        ((soc1.lsu.io_core_exe_0_req_bits_uop_uses_stq == 1'b1)
                        ?
                          (
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h0 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_0_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h1 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_1_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h2 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_2_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h3 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_3_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h4 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_4_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h5 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_5_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h6 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_6_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h7 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_7_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h8 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_8_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h9 ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_9_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'ha ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_10_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'hb ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_11_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'hc ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_12_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'hd ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_13_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'he ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_14_bits_uop_rob_idx) : 1'b1) &&
                          (soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'hf ? !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_15_bits_uop_rob_idx) : 1'b1)
                          )
                        :
                        1'b1)

                      : 1'b1;


	wire ME_4_lsufence;
	assign ME_4_lsufence = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
                      soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx == soc2.lsu.io_core_exe_0_req_bits_uop_rob_idx &&
										( soc1.lsu.io_core_exe_0_req_bits_sfence_bits_addr != soc2.lsu.io_core_exe_0_req_bits_sfence_bits_addr ||
											soc1.lsu.io_core_exe_0_req_bits_sfence_bits_rs1 != soc2.lsu.io_core_exe_0_req_bits_sfence_bits_rs1 ||
											soc1.lsu.io_core_exe_0_req_bits_sfence_bits_rs2 != soc2.lsu.io_core_exe_0_req_bits_sfence_bits_rs2 ) ) ?
											isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx) == 1'b0 : 1'b1;


	wire ME_4_lsufp;
	assign ME_4_lsufp = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
                        soc1.lsu.io_core_fp_stdata_bits_uop_rob_idx == soc2.lsu.io_core_fp_stdata_bits_uop_rob_idx &&
											( soc1.lsu.io_core_fp_stdata_bits_data != soc2.lsu.io_core_fp_stdata_bits_data) ) ?
											isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.io_core_fp_stdata_bits_uop_rob_idx) == 1'b0 : 1'b1;

  wire ME_4_lcam_st;
  assign ME_4_lcam_st = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
                        (soc1.lsu.do_st_search_0 == 1'b1) && (soc2.lsu.do_st_search_0 == 1'b1) && (soc1.lsu.lcam_stq_idx_0 == soc2.lsu.lcam_stq_idx_0) &&
                      ( soc1.lsu.lcam_addr_0 != soc2.lsu.lcam_addr_0) ) ?
                      isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.lsu.lcam_stq_idx_0]) == 1'b0 : 1'b1;

  wire ME_4_lcam_ld;
  assign ME_4_lcam_ld = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
                        (soc1.lsu.do_ld_search_0 == 1'b1) && (soc2.lsu.do_ld_search_0 == 1'b1) && (soc1.lsu.lcam_ldq_idx_0 == soc2.lsu.lcam_ldq_idx_0) &&
                      ( soc1.lsu.lcam_addr_0 != soc2.lsu.lcam_addr_0) ) ?
                      isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.lsu.lcam_ldq_idx_0]) == 1'b0 : 1'b1;
                      
      wire ME_4_lsu_iresp;
      assign ME_4_lsu_iresp = /*((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && !root_id_killed && !root_id_already_killed) &&*/
      				soc1.lsu.io_core_exe_0_iresp_bits_uop_rob_idx == soc2.lsu.io_core_exe_0_iresp_bits_uop_rob_idx &&
      				soc1.lsu.io_core_exe_0_iresp_bits_data != soc2.lsu.io_core_exe_0_iresp_bits_data
      				?
      					!isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.io_core_exe_0_iresp_bits_uop_rob_idx)
      				:
      				1'b1;
      				
      wire ME_4_MemAddrCalc;
      assign ME_4_MemAddrCalc = /*((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && !root_id_killed && !root_id_already_killed) &&*/
      				soc1.core.mem_units_0.maddrcalc.io_req_bits_uop_rob_idx == soc2.core.mem_units_0.maddrcalc.io_req_bits_uop_rob_idx &&
      				(soc1.core.mem_units_0.maddrcalc.io_req_bits_rs1_data != soc2.core.mem_units_0.maddrcalc.io_req_bits_rs1_data ||
      				soc1.core.mem_units_0.maddrcalc.io_req_bits_rs2_data != soc2.core.mem_units_0.maddrcalc.io_req_bits_rs2_data)
      				?
      					!isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_units_0.maddrcalc.io_req_bits_uop_rob_idx)
      				:
      				1'b1;
      				
                      

	wire ME_4;
	assign ME_4 = ME_4_alu && ME_4_div && ME_4_fpiu && ME_4_jmpalu && ME_4_ifpu && ME_4_imul && ME_4_lsu && ME_4_lsufence && ME_4_lsufp & ME_4_lcam_st & ME_4_lcam_ld & ME_4_lsu_iresp & ME_4_MemAddrCalc;
	
	wire ME_4_new_alu;
	assign ME_4_new_alu = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	soc1.core.csr_exe_unit.alu.io_req_bits_uop_rob_idx == soc2.core.csr_exe_unit.alu.io_req_bits_uop_rob_idx &&
	(  soc1.core.csr_exe_unit.alu.io_req_bits_rs1_data != soc2.core.csr_exe_unit.alu.io_req_bits_rs1_data ||
		soc1.core.csr_exe_unit.alu.io_req_bits_rs2_data != soc2.core.csr_exe_unit.alu.io_req_bits_rs2_data ) ) ?
		!ROBisOlder(soc1.core.csr_exe_unit.alu.io_req_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.core.csr_exe_unit.alu.io_req_bits_uop_rob_idx != root_id
		: 1'b1;
		
	wire ME_4_new_div;
	assign ME_4_new_div = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) && */
	soc1.core.csr_exe_unit.div.io_req_bits_uop_rob_idx == soc2.core.csr_exe_unit.div.io_req_bits_uop_rob_idx &&
	( soc1.core.csr_exe_unit.div.io_req_bits_rs1_data != soc2.core.csr_exe_unit.div.io_req_bits_rs1_data ||
		soc1.core.csr_exe_unit.div.io_req_bits_rs2_data != soc2.core.csr_exe_unit.div.io_req_bits_rs2_data ) ) ?
		!ROBisOlder(soc1.core.csr_exe_unit.div.io_req_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.core.csr_exe_unit.div.io_req_bits_uop_rob_idx != root_id &&
		!ROBisOlder(soc1.core.csr_exe_unit.div.io_req_bits_uop_yrot, root_id,soc1.core.rob.io_rob_head_idx) && soc1.core.csr_exe_unit.div.io_req_bits_uop_yrot != root_id
		: 1'b1;
			
			
	wire ME_4_new_fpiu;
	assign ME_4_new_fpiu =  (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	soc1.core.fp_pipeline.fpiu_unit.io_req_bits_uop_rob_idx == soc2.core.fp_pipeline.fpiu_unit.io_req_bits_uop_rob_idx &&
	( soc1.core.fp_pipeline.fpiu_unit.io_req_bits_rs1_data != soc2.core.fp_pipeline.fpiu_unit.io_req_bits_rs1_data ||
		soc1.core.fp_pipeline.fpiu_unit.io_req_bits_rs2_data != soc2.core.fp_pipeline.fpiu_unit.io_req_bits_rs2_data ||
		soc1.core.fp_pipeline.fpiu_unit.io_req_bits_rs3_data != soc2.core.fp_pipeline.fpiu_unit.io_req_bits_rs3_data ) ) ?
		!ROBisOlder(soc1.core.fp_pipeline.fpiu_unit.io_req_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.core.fp_pipeline.fpiu_unit.io_req_bits_uop_rob_idx != root_id
		: 1'b1;
				
				
	wire ME_4_new_jmpalu;
	assign ME_4_new_jmpalu =  (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	soc1.core.jmp_unit.alu.io_req_bits_uop_rob_idx == soc2.core.jmp_unit.alu.io_req_bits_uop_rob_idx &&
	( soc1.core.jmp_unit.alu.io_req_bits_rs1_data != soc2.core.jmp_unit.alu.io_req_bits_rs1_data ||
		soc1.core.jmp_unit.alu.io_req_bits_rs2_data != soc2.core.jmp_unit.alu.io_req_bits_rs2_data ) ) ?
		!ROBisOlder(soc1.core.jmp_unit.alu.io_req_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.core.jmp_unit.alu.io_req_bits_uop_rob_idx != root_id &&
		!ROBisOlder(soc1.core.jmp_unit.alu.io_req_bits_uop_yrot, root_id,soc1.core.rob.io_rob_head_idx) && soc1.core.jmp_unit.alu.io_req_bits_uop_yrot != root_id
		: 1'b1;
					
					
	wire ME_4_new_ifpu;
	assign ME_4_new_ifpu =  (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	soc1.core.jmp_unit.ifpu.io_req_bits_uop_rob_idx == soc2.core.jmp_unit.ifpu.io_req_bits_uop_rob_idx &&
	( soc1.core.jmp_unit.ifpu.io_req_bits_rs1_data != soc2.core.jmp_unit.ifpu.io_req_bits_rs1_data ) ) ?
	!ROBisOlder(soc1.core.jmp_unit.ifpu.io_req_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.core.jmp_unit.ifpu.io_req_bits_uop_rob_idx != root_id
	: 1'b1;


	wire ME_4_new_imul;
	assign ME_4_new_imul =  (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	soc1.core.jmp_unit.imul.io_req_bits_uop_rob_idx == soc2.core.jmp_unit.imul.io_req_bits_uop_rob_idx &&
	( soc1.core.jmp_unit.imul.io_req_bits_rs1_data != soc2.core.jmp_unit.imul.io_req_bits_rs1_data ||
		soc1.core.jmp_unit.imul.io_req_bits_rs2_data != soc2.core.jmp_unit.imul.io_req_bits_rs2_data ) ) ?
		!ROBisOlder(soc1.core.jmp_unit.imul.io_req_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.core.jmp_unit.imul.io_req_bits_uop_rob_idx != root_id
		: 1'b1;
		
		
	wire ME_4_new_lsu;
	assign ME_4_new_lsu = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx == soc2.lsu.io_core_exe_0_req_bits_uop_rob_idx &&
	( soc1.lsu.io_core_exe_0_req_bits_addr != soc2.lsu.io_core_exe_0_req_bits_addr ||
		soc1.lsu.io_core_exe_0_req_bits_data != soc2.lsu.io_core_exe_0_req_bits_data ) )
		?
		!ROBisOlder(soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx != root_id &&
		
		((soc1.lsu.io_core_exe_0_req_bits_uop_uses_ldq == 1'b1)
		?
		(
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h0 ? !ROBisOlder(soc1.lsu.ldq_0_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_0_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h1 ? !ROBisOlder(soc1.lsu.ldq_1_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_1_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h2 ? !ROBisOlder(soc1.lsu.ldq_2_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_2_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h3 ? !ROBisOlder(soc1.lsu.ldq_3_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_3_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h4 ? !ROBisOlder(soc1.lsu.ldq_4_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_4_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h5 ? !ROBisOlder(soc1.lsu.ldq_5_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_5_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h6 ? !ROBisOlder(soc1.lsu.ldq_6_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_6_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h7 ? !ROBisOlder(soc1.lsu.ldq_7_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_7_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h8 ? !ROBisOlder(soc1.lsu.ldq_8_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_8_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'h9 ? !ROBisOlder(soc1.lsu.ldq_9_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_9_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'hb ? !ROBisOlder(soc1.lsu.ldq_10_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_10_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'ha ? !ROBisOlder(soc1.lsu.ldq_11_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_11_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'hc ? !ROBisOlder(soc1.lsu.ldq_12_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_12_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'hd ? !ROBisOlder(soc1.lsu.ldq_13_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_13_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'he ? !ROBisOlder(soc1.lsu.ldq_14_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_14_bits_uop_rob_idx != root_id : 1'b1) &&
			(soc1.lsu.io_core_exe_0_req_bits_uop_ldq_idx == 4'hf ? !ROBisOlder(soc1.lsu.ldq_15_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.ldq_15_bits_uop_rob_idx != root_id : 1'b1)
			)
			:
			1'b1)&&
			
			((soc1.lsu.io_core_exe_0_req_bits_uop_uses_stq == 1'b1)
			?
			(
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h0 ? !ROBisOlder(soc1.lsu.stq_0_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_0_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h1 ? !ROBisOlder(soc1.lsu.stq_1_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_1_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h2 ? !ROBisOlder(soc1.lsu.stq_2_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_2_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h3 ? !ROBisOlder(soc1.lsu.stq_3_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_3_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h4 ? !ROBisOlder(soc1.lsu.stq_4_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_4_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h5 ? !ROBisOlder(soc1.lsu.stq_5_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_5_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h6 ? !ROBisOlder(soc1.lsu.stq_6_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_6_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h7 ? !ROBisOlder(soc1.lsu.stq_7_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_7_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h8 ? !ROBisOlder(soc1.lsu.stq_8_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_8_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'h9 ? !ROBisOlder(soc1.lsu.stq_9_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_9_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'ha ? !ROBisOlder(soc1.lsu.stq_10_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_10_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'hb ? !ROBisOlder(soc1.lsu.stq_11_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_11_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'hc ? !ROBisOlder(soc1.lsu.stq_12_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_12_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'hd ? !ROBisOlder(soc1.lsu.stq_13_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_13_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'he ? !ROBisOlder(soc1.lsu.stq_14_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_14_bits_uop_rob_idx != root_id : 1'b1) &&
				(soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx == 4'hf ? !ROBisOlder(soc1.lsu.stq_15_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.stq_15_bits_uop_rob_idx != root_id : 1'b1)
				)
				:
				1'b1)
				
				: 1'b1;
					
					
	wire ME_4_new_lsufence;
	assign ME_4_new_lsufence = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx == soc2.lsu.io_core_exe_0_req_bits_uop_rob_idx &&
	( soc1.lsu.io_core_exe_0_req_bits_sfence_bits_addr != soc2.lsu.io_core_exe_0_req_bits_sfence_bits_addr ||
		soc1.lsu.io_core_exe_0_req_bits_sfence_bits_rs1 != soc2.lsu.io_core_exe_0_req_bits_sfence_bits_rs1 ||
		soc1.lsu.io_core_exe_0_req_bits_sfence_bits_rs2 != soc2.lsu.io_core_exe_0_req_bits_sfence_bits_rs2 ) ) ?
		!ROBisOlder(soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.io_core_exe_0_req_bits_uop_rob_idx != root_id 
		: 1'b1;
						
						
	wire ME_4_new_lsufp;
	assign ME_4_new_lsufp = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	soc1.lsu.io_core_fp_stdata_bits_uop_rob_idx == soc2.lsu.io_core_fp_stdata_bits_uop_rob_idx &&
	( soc1.lsu.io_core_fp_stdata_bits_data != soc2.lsu.io_core_fp_stdata_bits_data) ) ?
	!ROBisOlder(soc1.lsu.io_core_fp_stdata_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.io_core_fp_stdata_bits_uop_rob_idx != root_id 
	: 1'b1;

	wire ME_4_new_lcam_st;
	assign ME_4_new_lcam_st = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	(soc1.lsu.do_st_search_0 == 1'b1) && (soc2.lsu.do_st_search_0 == 1'b1) && (soc1.lsu.lcam_stq_idx_0 == soc2.lsu.lcam_stq_idx_0) &&
	( soc1.lsu.lcam_addr_0 != soc2.lsu.lcam_addr_0) ) ?
	!ROBisOlder(stq_rob_idx_1[soc1.lsu.lcam_stq_idx_0], root_id,soc1.core.rob.io_rob_head_idx) && stq_rob_idx_1[soc1.lsu.lcam_stq_idx_0] != root_id 

	: 1'b1;

	wire ME_4_new_lcam_ld;
	assign ME_4_new_lcam_ld = (/* ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed)) &&*/
	(soc1.lsu.do_ld_search_0 == 1'b1) && (soc2.lsu.do_ld_search_0 == 1'b1) && (soc1.lsu.lcam_ldq_idx_0 == soc2.lsu.lcam_ldq_idx_0) &&
	( soc1.lsu.lcam_addr_0 != soc2.lsu.lcam_addr_0) ) ?
	!ROBisOlder(ldq_rob_idx_1[soc1.lsu.lcam_ldq_idx_0], root_id,soc1.core.rob.io_rob_head_idx) && ldq_rob_idx_1[soc1.lsu.lcam_ldq_idx_0] != root_id 
	: 1'b1;

	wire ME_4_new_lsu_iresp;
	assign ME_4_new_lsu_iresp = /*((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && !root_id_killed && !root_id_already_killed) &&*/
	soc1.lsu.io_core_exe_0_iresp_bits_uop_rob_idx == soc2.lsu.io_core_exe_0_iresp_bits_uop_rob_idx &&
	soc1.lsu.io_core_exe_0_iresp_bits_data != soc2.lsu.io_core_exe_0_iresp_bits_data
	?
	!ROBisOlder(soc1.lsu.io_core_exe_0_iresp_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.lsu.io_core_exe_0_iresp_bits_uop_rob_idx != root_id 
	:
	1'b1;

	wire ME_4_new_MemAddrCalc;
	assign ME_4_new_MemAddrCalc = /*((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && !root_id_killed && !root_id_already_killed) &&*/
	soc1.core.mem_units_0.maddrcalc.io_req_bits_uop_rob_idx == soc2.core.mem_units_0.maddrcalc.io_req_bits_uop_rob_idx &&
	(soc1.core.mem_units_0.maddrcalc.io_req_bits_rs1_data != soc2.core.mem_units_0.maddrcalc.io_req_bits_rs1_data ||
		soc1.core.mem_units_0.maddrcalc.io_req_bits_rs2_data != soc2.core.mem_units_0.maddrcalc.io_req_bits_rs2_data)
		?
		!ROBisOlder(soc1.core.mem_units_0.maddrcalc.io_req_bits_uop_rob_idx, root_id,soc1.core.rob.io_rob_head_idx) && soc1.core.mem_units_0.maddrcalc.io_req_bits_uop_rob_idx != root_id 
		:
		1'b1;
		
	wire ME_4_new;
	assign ME_4_new = ME_4_new_alu && ME_4_new_div && ME_4_new_fpiu && ME_4_new_jmpalu && ME_4_new_ifpu && ME_4_new_imul && ME_4_new_lsu && ME_4_new_lsufence && ME_4_new_lsufp & ME_4_new_lcam_st & ME_4_new_lcam_ld & ME_4_new_lsu_iresp & ME_4_new_MemAddrCalc;

//*******************************************//
//************ME-5 & ME-6********************//
//write one combinational process for both ME-5 and ME-6
//for every ROB slot or bookkeeping buffer:
//check if stored ROB ID is committable
//store branch mask in corresponding variable
//set the other variable to default value (12'hfff for uncommitable tags, 12'h0 for committable tags)

//Soc1

  wire [11:0] alu_T_2_com_1;
  wire [11:0] alu_T_2_uncom_1;

  always @(*)
  begin
    alu_T_2_com_1 = 12'h0;
    alu_T_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.csr_exe_unit.alu.r_uops_0_rob_idx) && soc1.core.csr_exe_unit.alu.r_valids_0)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.csr_exe_unit.alu.r_uops_0_rob_idx))
      begin
        alu_T_2_com_1 = soc1.core.csr_exe_unit.alu.r_uops_0_br_mask;
        alu_T_2_uncom_1 = 12'hfff;
      end
      else
      begin
        alu_T_2_com_1 = 12'h0;
        alu_T_2_uncom_1 = soc1.core.csr_exe_unit.alu.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] div_r_com_1;
  wire [11:0] div_r_uncom_1;

  always @(*)
  begin
    div_r_com_1 = 12'h0;
    div_r_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.csr_exe_unit.div.r_uop_rob_idx) && (soc1.core.csr_exe_unit.div.div.state == 3'h3))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.csr_exe_unit.div.r_uop_rob_idx))
      begin
        div_r_com_1 = soc1.core.csr_exe_unit.div.r_uop_br_mask;
        div_r_uncom_1 = 12'hfff;
      end
      else
      begin
        div_r_com_1 = 12'h0;
        div_r_uncom_1 = soc1.core.csr_exe_unit.div.r_uop_br_mask;
      end
    end
  end

  wire [11:0] exe_reg_0_com_1;
  wire [11:0] exe_reg_0_uncom_1;

  always @(*)
  begin
    exe_reg_0_com_1 = 12'h0;
    exe_reg_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.iregister_read.exe_reg_uops_0_rob_idx) && soc1.core.iregister_read.exe_reg_valids_0 && !(soc1.core.iregister_read.exe_reg_uops_0_uses_stq && stq_committed_1[soc1.core.iregister_read.exe_reg_uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.exe_reg_uops_0_rob_idx))
      begin
        exe_reg_0_com_1 = soc1.core.iregister_read.exe_reg_uops_0_br_mask;
        exe_reg_0_uncom_1 = 12'hfff;
      end
      else
      begin
        exe_reg_0_com_1 = 12'h0;
        exe_reg_0_uncom_1 = soc1.core.iregister_read.exe_reg_uops_0_br_mask;
      end
    end
  end

  wire [11:0] exe_reg_1_com_1;
  wire [11:0] exe_reg_1_uncom_1;

  always @(*)
  begin
    exe_reg_1_com_1 = 12'h0;
    exe_reg_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.iregister_read.exe_reg_uops_1_rob_idx) && soc1.core.iregister_read.exe_reg_valids_1 && !(soc1.core.iregister_read.exe_reg_uops_1_uses_stq && stq_committed_1[soc1.core.iregister_read.exe_reg_uops_1_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.exe_reg_uops_1_rob_idx))
      begin
        exe_reg_1_com_1 = soc1.core.iregister_read.exe_reg_uops_1_br_mask;
        exe_reg_1_uncom_1 = 12'hfff;
      end
      else
      begin
        exe_reg_1_com_1 = 12'h0;
        exe_reg_1_uncom_1 = soc1.core.iregister_read.exe_reg_uops_1_br_mask;
      end
    end
  end

  wire [11:0] exe_reg_2_com_1;
  wire [11:0] exe_reg_2_uncom_1;

  always @(*)
  begin
    exe_reg_2_com_1 = 12'h0;
    exe_reg_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.iregister_read.exe_reg_uops_2_rob_idx) && soc1.core.iregister_read.exe_reg_valids_2 && !(soc1.core.iregister_read.exe_reg_uops_2_uses_stq && stq_committed_1[soc1.core.iregister_read.exe_reg_uops_2_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.exe_reg_uops_2_rob_idx))
      begin
        exe_reg_2_com_1 = soc1.core.iregister_read.exe_reg_uops_2_br_mask;
        exe_reg_2_uncom_1 = 12'hfff;
      end
      else
      begin
        exe_reg_2_com_1 = 12'h0;
        exe_reg_2_uncom_1 = soc1.core.iregister_read.exe_reg_uops_2_br_mask;
      end
    end
  end

  wire [11:0] rrd_0_com_1;
  wire [11:0] rrd_0_uncom_1;

  always @(*)
  begin
    rrd_0_com_1 = 12'h0;
    rrd_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.iregister_read.rrd_uops_0_REG_rob_idx) && soc1.core.iregister_read.rrd_valids_0_REG && !(soc1.core.iregister_read.rrd_uops_0_REG_uses_stq && stq_committed_1[soc1.core.iregister_read.rrd_uops_0_REG_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.rrd_uops_0_REG_rob_idx))
      begin
        rrd_0_com_1 = soc1.core.iregister_read.rrd_uops_0_REG_br_mask;
        rrd_0_uncom_1 = 12'hfff;
      end
      else
      begin
        rrd_0_com_1 = 12'h0;
        rrd_0_uncom_1 = soc1.core.iregister_read.rrd_uops_0_REG_br_mask;
      end
    end
  end

  wire [11:0] rrd_1_com_1;
  wire [11:0] rrd_1_uncom_1;

  always @(*)
  begin
    rrd_1_com_1 = 12'h0;
    rrd_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.iregister_read.rrd_uops_1_REG_rob_idx) && soc1.core.iregister_read.rrd_valids_1_REG && !(soc1.core.iregister_read.rrd_uops_1_REG_uses_stq && stq_committed_1[soc1.core.iregister_read.rrd_uops_1_REG_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.rrd_uops_1_REG_rob_idx))
      begin
        rrd_1_com_1 = soc1.core.iregister_read.rrd_uops_1_REG_br_mask;
        rrd_1_uncom_1 = 12'hfff;
      end
      else
      begin
        rrd_1_com_1 = 12'h0;
        rrd_1_uncom_1 = soc1.core.iregister_read.rrd_uops_1_REG_br_mask;
      end
    end
  end

  wire [11:0] rrd_2_com_1;
  wire [11:0] rrd_2_uncom_1;

  always @(*)
  begin
    rrd_2_com_1 = 12'h0;
    rrd_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.iregister_read.rrd_uops_2_REG_rob_idx) && soc1.core.iregister_read.rrd_valids_2_REG && !(soc1.core.iregister_read.rrd_uops_2_REG_uses_stq && stq_committed_1[soc1.core.iregister_read.rrd_uops_2_REG_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.rrd_uops_2_REG_rob_idx))
      begin
        rrd_2_com_1 = soc1.core.iregister_read.rrd_uops_2_REG_br_mask;
        rrd_2_uncom_1 = 12'hfff;
      end
      else
      begin
        rrd_2_com_1 = 12'h0;
        rrd_2_uncom_1 = soc1.core.iregister_read.rrd_uops_2_REG_br_mask;
      end
    end
  end

  wire [11:0] bkq_0_com_1;
  wire [11:0] bkq_0_uncom_1;

  always @(*)
  begin
    bkq_0_com_1 = 12'h0;
    bkq_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.queue.uops_0_rob_idx) && soc1.core.jmp_unit.queue.valids_0 /*&& !(soc1.core.jmp_unit.queue.uops_0_uses_stq && stq_committed_1[soc1.core.jmp_unit.queue.uops_0_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.queue.uops_0_rob_idx))
      begin
        bkq_0_com_1 = soc1.core.jmp_unit.queue.uops_0_br_mask;
        bkq_0_uncom_1 = 12'hfff;
      end
      else
      begin
        bkq_0_com_1 = 12'h0;
        bkq_0_uncom_1 = soc1.core.jmp_unit.queue.uops_0_br_mask;
      end
    end
  end

  wire [11:0] bkq_1_com_1;
  wire [11:0] bkq_1_uncom_1;

  always @(*)
  begin
    bkq_1_com_1 = 12'h0;
    bkq_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.queue.uops_1_rob_idx) && soc1.core.jmp_unit.queue.valids_1 /*&& !(soc1.core.jmp_unit.queue.uops_1_uses_stq && stq_committed_1[soc1.core.jmp_unit.queue.uops_1_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.queue.uops_1_rob_idx))
      begin
        bkq_1_com_1 = soc1.core.jmp_unit.queue.uops_1_br_mask;
        bkq_1_uncom_1 = 12'hfff;
      end
      else
      begin
        bkq_1_com_1 = 12'h0;
        bkq_1_uncom_1 = soc1.core.jmp_unit.queue.uops_1_br_mask;
      end
    end
  end

  wire [11:0] bkq_2_com_1;
  wire [11:0] bkq_2_uncom_1;

  always @(*)
  begin
    bkq_2_com_1 = 12'h0;
    bkq_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.queue.uops_2_rob_idx) && soc1.core.jmp_unit.queue.valids_2 /*&& !(soc1.core.jmp_unit.queue.uops_2_uses_stq && stq_committed_1[soc1.core.jmp_unit.queue.uops_2_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.queue.uops_2_rob_idx))
      begin
        bkq_2_com_1 = soc1.core.jmp_unit.queue.uops_2_br_mask;
        bkq_2_uncom_1 = 12'hfff;
      end
      else
      begin
        bkq_2_com_1 = 12'h0;
        bkq_2_uncom_1 = soc1.core.jmp_unit.queue.uops_2_br_mask;
      end
    end
  end

  wire [11:0] bkq_3_com_1;
  wire [11:0] bkq_3_uncom_1;

  always @(*)
  begin
    bkq_3_com_1 = 12'h0;
    bkq_3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.queue.uops_3_rob_idx) && soc1.core.jmp_unit.queue.valids_3 /*&& !(soc1.core.jmp_unit.queue.uops_3_uses_stq && stq_committed_1[soc1.core.jmp_unit.queue.uops_3_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.queue.uops_3_rob_idx))
      begin
        bkq_3_com_1 = soc1.core.jmp_unit.queue.uops_3_br_mask;
        bkq_3_uncom_1 = 12'hfff;
      end
      else
      begin
        bkq_3_com_1 = 12'h0;
        bkq_3_uncom_1 = soc1.core.jmp_unit.queue.uops_3_br_mask;
      end
    end
  end

  wire [11:0] bkq_4_com_1;
  wire [11:0] bkq_4_uncom_1;

  always @(*)
  begin
    bkq_4_com_1 = 12'h0;
    bkq_4_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.queue.uops_4_rob_idx) && soc1.core.jmp_unit.queue.valids_4 /*&& !(soc1.core.jmp_unit.queue.uops_4_uses_stq && stq_committed_1[soc1.core.jmp_unit.queue.uops_4_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.queue.uops_4_rob_idx))
      begin
        bkq_4_com_1 = soc1.core.jmp_unit.queue.uops_4_br_mask;
        bkq_4_uncom_1 = 12'hfff;
      end
      else
      begin
        bkq_4_com_1 = 12'h0;
        bkq_4_uncom_1 = soc1.core.jmp_unit.queue.uops_4_br_mask;
      end
    end
  end

  wire [11:0] alu_T_2_0_com_1;
  wire [11:0] alu_T_2_0_uncom_1;

  always @(*)
  begin
    alu_T_2_0_com_1 = 12'h0;
    alu_T_2_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.alu.r_uops_0_rob_idx) && soc1.core.jmp_unit.alu.r_valids_0)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.alu.r_uops_0_rob_idx))
      begin
        alu_T_2_0_com_1 = soc1.core.jmp_unit.alu.r_uops_0_br_mask;
        alu_T_2_0_uncom_1 = 12'hfff;
      end
      else
      begin
        alu_T_2_0_com_1 = 12'h0;
        alu_T_2_0_uncom_1 = soc1.core.jmp_unit.alu.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] alu_T_2_1_com_1;
  wire [11:0] alu_T_2_1_uncom_1;

  always @(*)
  begin
    alu_T_2_1_com_1 = 12'h0;
    alu_T_2_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.alu.r_uops_1_rob_idx) && soc1.core.jmp_unit.alu.r_valids_1)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.alu.r_uops_1_rob_idx))
      begin
        alu_T_2_1_com_1 = soc1.core.jmp_unit.alu.r_uops_1_br_mask;
        alu_T_2_1_uncom_1 = 12'hfff;
      end
      else
      begin
        alu_T_2_1_com_1 = 12'h0;
        alu_T_2_1_uncom_1 = soc1.core.jmp_unit.alu.r_uops_1_br_mask;
      end
    end
  end

  wire [11:0] alu_T_2_2_com_1;
  wire [11:0] alu_T_2_2_uncom_1;

  always @(*)
  begin
    alu_T_2_2_com_1 = 12'h0;
    alu_T_2_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.alu.r_uops_2_rob_idx) && soc1.core.jmp_unit.alu.r_valids_2)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.alu.r_uops_2_rob_idx))
      begin
        alu_T_2_2_com_1 = soc1.core.jmp_unit.alu.r_uops_2_br_mask;
        alu_T_2_2_uncom_1 = 12'hfff;
      end
      else
      begin
        alu_T_2_2_com_1 = 12'h0;
        alu_T_2_2_uncom_1 = soc1.core.jmp_unit.alu.r_uops_2_br_mask;
      end
    end
  end

  wire [11:0] ifpu_T_2_0_com_1;
  wire [11:0] ifpu_T_2_0_uncom_1;

  always @(*)
  begin
    ifpu_T_2_0_com_1 = 12'h0;
    ifpu_T_2_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.ifpu.r_uops_0_rob_idx) && soc1.core.jmp_unit.ifpu.r_valids_0 /*&& !(soc1.core.jmp_unit.ifpu.r_uops_0_uses_stq && stq_committed_1[soc1.core.jmp_unit.ifpu.r_uops_0_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.ifpu.r_uops_0_rob_idx))
      begin
        ifpu_T_2_0_com_1 = soc1.core.jmp_unit.ifpu.r_uops_0_br_mask;
        ifpu_T_2_0_uncom_1 = 12'hfff;
      end
      else
      begin
        ifpu_T_2_0_com_1 = 12'h0;
        ifpu_T_2_0_uncom_1 = soc1.core.jmp_unit.ifpu.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] ifpu_T_2_1_com_1;
  wire [11:0] ifpu_T_2_1_uncom_1;

  always @(*)
  begin
    ifpu_T_2_1_com_1 = 12'h0;
    ifpu_T_2_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.ifpu.r_uops_1_rob_idx) && soc1.core.jmp_unit.ifpu.r_valids_1 /*&& !(soc1.core.jmp_unit.ifpu.r_uops_1_uses_stq && stq_committed_1[soc1.core.jmp_unit.ifpu.r_uops_1_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.ifpu.r_uops_1_rob_idx))
      begin
        ifpu_T_2_1_com_1 = soc1.core.jmp_unit.ifpu.r_uops_1_br_mask;
        ifpu_T_2_1_uncom_1 = 12'hfff;
      end
      else
      begin
        ifpu_T_2_1_com_1 = 12'h0;
        ifpu_T_2_1_uncom_1 = soc1.core.jmp_unit.ifpu.r_uops_1_br_mask;
      end
    end
  end



  wire [11:0] imul_T_2_0_com_1;
  wire [11:0] imul_T_2_0_uncom_1;

  always @(*)
  begin
    imul_T_2_0_com_1 = 12'h0;
    imul_T_2_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.imul.r_uops_0_rob_idx) && soc1.core.jmp_unit.imul.r_valids_0)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.imul.r_uops_0_rob_idx))
      begin
        imul_T_2_0_com_1 = soc1.core.jmp_unit.imul.r_uops_0_br_mask;
        imul_T_2_0_uncom_1 = 12'hfff;
      end
      else
      begin
        imul_T_2_0_com_1 = 12'h0;
        imul_T_2_0_uncom_1 = soc1.core.jmp_unit.imul.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] imul_T_2_1_com_1;
  wire [11:0] imul_T_2_1_uncom_1;

  always @(*)
  begin
    imul_T_2_1_com_1 = 12'h0;
    imul_T_2_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.imul.r_uops_1_rob_idx) && soc1.core.jmp_unit.imul.r_valids_1)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.imul.r_uops_1_rob_idx))
      begin
        imul_T_2_1_com_1 = soc1.core.jmp_unit.imul.r_uops_1_br_mask;
        imul_T_2_1_uncom_1 = 12'hfff;
      end
      else
      begin
        imul_T_2_1_com_1 = 12'h0;
        imul_T_2_1_uncom_1 = soc1.core.jmp_unit.imul.r_uops_1_br_mask;
      end
    end
  end

  wire [11:0] imul_T_2_2_com_1;
  wire [11:0] imul_T_2_2_uncom_1;

  always @(*)
  begin
    imul_T_2_2_com_1 = 12'h0;
    imul_T_2_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.jmp_unit.imul.r_uops_2_rob_idx) && soc1.core.jmp_unit.imul.r_valids_2)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.imul.r_uops_2_rob_idx))
      begin
        imul_T_2_2_com_1 = soc1.core.jmp_unit.imul.r_uops_2_br_mask;
        imul_T_2_2_uncom_1 = 12'hfff;
      end
      else
      begin
        imul_T_2_2_com_1 = 12'h0;
        imul_T_2_2_uncom_1 = soc1.core.jmp_unit.imul.r_uops_2_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_0_com_1;
  wire [11:0] fp_issue_slot_0_uncom_1;

  always @(*)
  begin
    fp_issue_slot_0_com_1 = 12'h0;
    fp_issue_slot_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_0.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx))
      begin
        fp_issue_slot_0_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_br_mask;
        fp_issue_slot_0_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_0_com_1 = 12'h0;
        fp_issue_slot_0_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_1_com_1;
  wire [11:0] fp_issue_slot_1_uncom_1;

  always @(*)
  begin
    fp_issue_slot_1_com_1 = 12'h0;
    fp_issue_slot_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_1.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx))
      begin
        fp_issue_slot_1_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_br_mask;
        fp_issue_slot_1_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_1_com_1 = 12'h0;
        fp_issue_slot_1_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_2_com_1;
  wire [11:0] fp_issue_slot_2_uncom_1;

  always @(*)
  begin
    fp_issue_slot_2_com_1 = 12'h0;
    fp_issue_slot_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_2.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx))
      begin
        fp_issue_slot_2_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_br_mask;
        fp_issue_slot_2_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_2_com_1 = 12'h0;
        fp_issue_slot_2_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_3_com_1;
  wire [11:0] fp_issue_slot_3_uncom_1;

  always @(*)
  begin
    fp_issue_slot_3_com_1 = 12'h0;
    fp_issue_slot_3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_3.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx))
      begin
        fp_issue_slot_3_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_br_mask;
        fp_issue_slot_3_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_3_com_1 = 12'h0;
        fp_issue_slot_3_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_4_com_1;
  wire [11:0] fp_issue_slot_4_uncom_1;

  always @(*)
  begin
    fp_issue_slot_4_com_1 = 12'h0;
    fp_issue_slot_4_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_4.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx))
      begin
        fp_issue_slot_4_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_br_mask;
        fp_issue_slot_4_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_4_com_1 = 12'h0;
        fp_issue_slot_4_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_5_com_1;
  wire [11:0] fp_issue_slot_5_uncom_1;

  always @(*)
  begin
    fp_issue_slot_5_com_1 = 12'h0;
    fp_issue_slot_5_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_5.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx))
      begin
        fp_issue_slot_5_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_br_mask;
        fp_issue_slot_5_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_5_com_1 = 12'h0;
        fp_issue_slot_5_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_6_com_1;
  wire [11:0] fp_issue_slot_6_uncom_1;

  always @(*)
  begin
    fp_issue_slot_6_com_1 = 12'h0;
    fp_issue_slot_6_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_6.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx))
      begin
        fp_issue_slot_6_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_br_mask;
        fp_issue_slot_6_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_6_com_1 = 12'h0;
        fp_issue_slot_6_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_7_com_1;
  wire [11:0] fp_issue_slot_7_uncom_1;

  always @(*)
  begin
    fp_issue_slot_7_com_1 = 12'h0;
    fp_issue_slot_7_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_7.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx))
      begin
        fp_issue_slot_7_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_br_mask;
        fp_issue_slot_7_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_7_com_1 = 12'h0;
        fp_issue_slot_7_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_8_com_1;
  wire [11:0] fp_issue_slot_8_uncom_1;

  always @(*)
  begin
    fp_issue_slot_8_com_1 = 12'h0;
    fp_issue_slot_8_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_8.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx))
      begin
        fp_issue_slot_8_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_br_mask;
        fp_issue_slot_8_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_8_com_1 = 12'h0;
        fp_issue_slot_8_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_9_com_1;
  wire [11:0] fp_issue_slot_9_uncom_1;

  always @(*)
  begin
    fp_issue_slot_9_com_1 = 12'h0;
    fp_issue_slot_9_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_9.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx))
      begin
        fp_issue_slot_9_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_br_mask;
        fp_issue_slot_9_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_9_com_1 = 12'h0;
        fp_issue_slot_9_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_10_com_1;
  wire [11:0] fp_issue_slot_10_uncom_1;

  always @(*)
  begin
    fp_issue_slot_10_com_1 = 12'h0;
    fp_issue_slot_10_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_10.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx))
      begin
        fp_issue_slot_10_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_br_mask;
        fp_issue_slot_10_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_10_com_1 = 12'h0;
        fp_issue_slot_10_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_11_com_1;
  wire [11:0] fp_issue_slot_11_uncom_1;

  always @(*)
  begin
    fp_issue_slot_11_com_1 = 12'h0;
    fp_issue_slot_11_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_11.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx))
      begin
        fp_issue_slot_11_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_br_mask;
        fp_issue_slot_11_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_11_com_1 = 12'h0;
        fp_issue_slot_11_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_12_com_1;
  wire [11:0] fp_issue_slot_12_uncom_1;

  always @(*)
  begin
    fp_issue_slot_12_com_1 = 12'h0;
    fp_issue_slot_12_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_12.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx))
      begin
        fp_issue_slot_12_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_br_mask;
        fp_issue_slot_12_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_12_com_1 = 12'h0;
        fp_issue_slot_12_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_13_com_1;
  wire [11:0] fp_issue_slot_13_uncom_1;

  always @(*)
  begin
    fp_issue_slot_13_com_1 = 12'h0;
    fp_issue_slot_13_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_13.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx))
      begin
        fp_issue_slot_13_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_br_mask;
        fp_issue_slot_13_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_13_com_1 = 12'h0;
        fp_issue_slot_13_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_14_com_1;
  wire [11:0] fp_issue_slot_14_uncom_1;

  always @(*)
  begin
    fp_issue_slot_14_com_1 = 12'h0;
    fp_issue_slot_14_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_14.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx))
      begin
        fp_issue_slot_14_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_br_mask;
        fp_issue_slot_14_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_14_com_1 = 12'h0;
        fp_issue_slot_14_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_15_com_1;
  wire [11:0] fp_issue_slot_15_uncom_1;

  always @(*)
  begin
    fp_issue_slot_15_com_1 = 12'h0;
    fp_issue_slot_15_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx) && soc1.core.fp_pipeline.fp_issue_unit.slots_15.io_valid && !(soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx))
      begin
        fp_issue_slot_15_com_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_br_mask;
        fp_issue_slot_15_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_15_com_1 = 12'h0;
        fp_issue_slot_15_uncom_1 = soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_0_com_1;
  wire [11:0] fp_bkq_0_uncom_1;

  always @(*)
  begin
    fp_bkq_0_com_1 = 12'h0;
    fp_bkq_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.queue.valids_0 && !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx))
      begin
        fp_bkq_0_com_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_br_mask;
        fp_bkq_0_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_0_com_1 = 12'h0;
        fp_bkq_0_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_1_com_1;
  wire [11:0] fp_bkq_1_uncom_1;

  always @(*)
  begin
    fp_bkq_1_com_1 = 12'h0;
    fp_bkq_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.queue.valids_1 && !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx))
      begin
        fp_bkq_1_com_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_br_mask;
        fp_bkq_1_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_1_com_1 = 12'h0;
        fp_bkq_1_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_2_com_1;
  wire [11:0] fp_bkq_2_uncom_1;

  always @(*)
  begin
    fp_bkq_2_com_1 = 12'h0;
    fp_bkq_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.queue.valids_2 && !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx))
      begin
        fp_bkq_2_com_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_br_mask;
        fp_bkq_2_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_2_com_1 = 12'h0;
        fp_bkq_2_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_3_com_1;
  wire [11:0] fp_bkq_3_uncom_1;

  always @(*)
  begin
    fp_bkq_3_com_1 = 12'h0;
    fp_bkq_3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.queue.valids_3 && !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx))
      begin
        fp_bkq_3_com_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_br_mask;
        fp_bkq_3_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_3_com_1 = 12'h0;
        fp_bkq_3_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_4_com_1;
  wire [11:0] fp_bkq_4_uncom_1;

  always @(*)
  begin
    fp_bkq_4_com_1 = 12'h0;
    fp_bkq_4_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.queue.valids_4 && !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx))
      begin
        fp_bkq_4_com_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_br_mask;
        fp_bkq_4_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_4_com_1 = 12'h0;
        fp_bkq_4_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_5_com_1;
  wire [11:0] fp_bkq_5_uncom_1;

  always @(*)
  begin
    fp_bkq_5_com_1 = 12'h0;
    fp_bkq_5_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.queue.valids_5 && !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx))
      begin
        fp_bkq_5_com_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_br_mask;
        fp_bkq_5_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_5_com_1 = 12'h0;
        fp_bkq_5_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_6_com_1;
  wire [11:0] fp_bkq_6_uncom_1;

  always @(*)
  begin
    fp_bkq_6_com_1 = 12'h0;
    fp_bkq_6_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.queue.valids_6 && !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx))
      begin
        fp_bkq_6_com_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_br_mask;
        fp_bkq_6_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_6_com_1 = 12'h0;
        fp_bkq_6_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_1_0_com_1;
  wire [11:0] fp_bkq_1_0_uncom_1;

  always @(*)
  begin
    fp_bkq_1_0_com_1 = 12'h0;
    fp_bkq_1_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0 && !(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx))
      begin
        fp_bkq_1_0_com_1 = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_br_mask;
        fp_bkq_1_0_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_1_0_com_1 = 12'h0;
        fp_bkq_1_0_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_1_1_com_1;
  wire [11:0] fp_bkq_1_1_uncom_1;

  always @(*)
  begin
    fp_bkq_1_1_com_1 = 12'h0;
    fp_bkq_1_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx)  && soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1 && !(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx))
      begin
        fp_bkq_1_1_com_1 = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_br_mask;
        fp_bkq_1_1_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_1_1_com_1 = 12'h0;
        fp_bkq_1_1_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_1_2_com_1;
  wire [11:0] fp_bkq_1_2_uncom_1;

  always @(*)
  begin
    fp_bkq_1_2_com_1 = 12'h0;
    fp_bkq_1_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2 && !(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx))
      begin
        fp_bkq_1_2_com_1 = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_br_mask;
        fp_bkq_1_2_uncom_1 = 12'hfff;
      end
      else
      begin
        fp_bkq_1_2_com_1 = 12'h0;
        fp_bkq_1_2_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_br_mask;
      end
    end
  end

  wire [11:0] fdiv_buf_com_1;
  wire [11:0] fdiv_buf_uncom_1;

  always @(*)
  begin
    fdiv_buf_com_1 = 12'h0;
    fdiv_buf_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_val)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx))
      begin
        fdiv_buf_com_1 = soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_br_mask;
        fdiv_buf_uncom_1 = 12'hfff;
      end
      else
      begin
        fdiv_buf_com_1 = 12'h0;
        fdiv_buf_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_br_mask;
      end
    end
  end

  wire [11:0] fdiv_divsqrt_com_1;
  wire [11:0] fdiv_divsqrt_uncom_1;

  always @(*)
  begin
    fdiv_divsqrt_com_1 = 12'h0;
    fdiv_divsqrt_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx))
      begin
        fdiv_divsqrt_com_1 = soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_br_mask;
        fdiv_divsqrt_uncom_1 = 12'hfff;
      end
      else
      begin
        fdiv_divsqrt_com_1 = 12'h0;
        fdiv_divsqrt_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_br_mask;
      end
    end
  end

  wire [11:0] fdiv_out_com_1;
  wire [11:0] fdiv_out_uncom_1;

  always @(*)
  begin
    fdiv_out_com_1 = 12'h0;
    fdiv_out_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_val)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx))
      begin
        fdiv_out_com_1 = soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_br_mask;
        fdiv_out_uncom_1 = 12'hfff;
      end
      else
      begin
        fdiv_out_com_1 = 12'h0;
        fdiv_out_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_br_mask;
      end
    end
  end

  wire [11:0] fpu_T_2_0_com_1;
  wire [11:0] fpu_T_2_0_uncom_1;

  always @(*)
  begin
    fpu_T_2_0_com_1 = 12'h0;
    fpu_T_2_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_0 && !(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx))
      begin
        fpu_T_2_0_com_1 = soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_br_mask;
        fpu_T_2_0_uncom_1 = 12'hfff;
      end
      else
      begin
        fpu_T_2_0_com_1 = 12'h0;
        fpu_T_2_0_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] fpu_T_2_1_com_1;
  wire [11:0] fpu_T_2_1_uncom_1;

  always @(*)
  begin
    fpu_T_2_1_com_1 = 12'h0;
    fpu_T_2_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_1 && !(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx))
      begin
        fpu_T_2_1_com_1 = soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_br_mask;
        fpu_T_2_1_uncom_1 = 12'hfff;
      end
      else
      begin
        fpu_T_2_1_com_1 = 12'h0;
        fpu_T_2_1_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_br_mask;
      end
    end
  end

  wire [11:0] fpu_T_2_2_com_1;
  wire [11:0] fpu_T_2_2_uncom_1;

  always @(*)
  begin
    fpu_T_2_2_com_1 = 12'h0;
    fpu_T_2_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_2 && !(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx))
      begin
        fpu_T_2_2_com_1 = soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_br_mask;
        fpu_T_2_2_uncom_1 = 12'hfff;
      end
      else
      begin
        fpu_T_2_2_com_1 = 12'h0;
        fpu_T_2_2_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_br_mask;
      end
    end
  end

  wire [11:0] fpu_T_2_3_com_1;
  wire [11:0] fpu_T_2_3_uncom_1;

  always @(*)
  begin
    fpu_T_2_3_com_1 = 12'h0;
    fpu_T_2_3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx) && soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_3 && !(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx))
      begin
        fpu_T_2_3_com_1 = soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_br_mask;
        fpu_T_2_3_uncom_1 = 12'hfff;
      end
      else
      begin
        fpu_T_2_3_com_1 = 12'h0;
        fpu_T_2_3_uncom_1 = soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_br_mask;
      end
    end
  end

  wire [11:0] f_exe_reg_com_1;
  wire [11:0] f_exe_reg_uncom_1;

  always @(*)
  begin
    f_exe_reg_com_1 = 12'h0;
    f_exe_reg_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx) && soc1.core.fp_pipeline.fregister_read.exe_reg_valids_0 && !(soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx))
      begin
        f_exe_reg_com_1 = soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_br_mask;
        f_exe_reg_uncom_1 = 12'hfff;
      end
      else
      begin
        f_exe_reg_com_1 = 12'h0;
        f_exe_reg_uncom_1 = soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_br_mask;
      end
    end
  end

  wire [11:0] f_rrd_com_1;
  wire [11:0] f_rrd_uncom_1;

  always @(*)
  begin
    f_rrd_com_1 = 12'h0;
    f_rrd_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx) && soc1.core.fp_pipeline.fregister_read.rrd_valids_0_REG && !(soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx))
      begin
        f_rrd_com_1 = soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_br_mask;
        f_rrd_uncom_1 = 12'hfff;
      end
      else
      begin
        f_rrd_com_1 = 12'h0;
        f_rrd_uncom_1 = soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_0_com_1;
  wire [11:0] int_issue_slot_0_uncom_1;

  always @(*)
  begin
    int_issue_slot_0_com_1 = 12'h0;
    int_issue_slot_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_0.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_0.io_valid && !(soc1.core.int_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_0.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_0.slot_uop_rob_idx))
      begin
        int_issue_slot_0_com_1 = soc1.core.int_issue_unit.slots_0.slot_uop_br_mask;
        int_issue_slot_0_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_0_com_1 = 12'h0;
        int_issue_slot_0_uncom_1 = soc1.core.int_issue_unit.slots_0.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_1_com_1;
  wire [11:0] int_issue_slot_1_uncom_1;

  always @(*)
  begin
    int_issue_slot_1_com_1 = 12'h0;
    int_issue_slot_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_1.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_1.io_valid && !(soc1.core.int_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_1.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_1.slot_uop_rob_idx))
      begin
        int_issue_slot_1_com_1 = soc1.core.int_issue_unit.slots_1.slot_uop_br_mask;
        int_issue_slot_1_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_1_com_1 = 12'h0;
        int_issue_slot_1_uncom_1 = soc1.core.int_issue_unit.slots_1.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_2_com_1;
  wire [11:0] int_issue_slot_2_uncom_1;

  always @(*)
  begin
    int_issue_slot_2_com_1 = 12'h0;
    int_issue_slot_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_2.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_2.io_valid && !(soc1.core.int_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_2.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_2.slot_uop_rob_idx))
      begin
        int_issue_slot_2_com_1 = soc1.core.int_issue_unit.slots_2.slot_uop_br_mask;
        int_issue_slot_2_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_2_com_1 = 12'h0;
        int_issue_slot_2_uncom_1 = soc1.core.int_issue_unit.slots_2.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_3_com_1;
  wire [11:0] int_issue_slot_3_uncom_1;

  always @(*)
  begin
    int_issue_slot_3_com_1 = 12'h0;
    int_issue_slot_3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_3.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_3.io_valid && !(soc1.core.int_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_3.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_3.slot_uop_rob_idx))
      begin
        int_issue_slot_3_com_1 = soc1.core.int_issue_unit.slots_3.slot_uop_br_mask;
        int_issue_slot_3_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_3_com_1 = 12'h0;
        int_issue_slot_3_uncom_1 = soc1.core.int_issue_unit.slots_3.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_4_com_1;
  wire [11:0] int_issue_slot_4_uncom_1;

  always @(*)
  begin
    int_issue_slot_4_com_1 = 12'h0;
    int_issue_slot_4_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_4.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_4.io_valid && !(soc1.core.int_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_4.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_4.slot_uop_rob_idx))
      begin
        int_issue_slot_4_com_1 = soc1.core.int_issue_unit.slots_4.slot_uop_br_mask;
        int_issue_slot_4_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_4_com_1 = 12'h0;
        int_issue_slot_4_uncom_1 = soc1.core.int_issue_unit.slots_4.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_5_com_1;
  wire [11:0] int_issue_slot_5_uncom_1;

  always @(*)
  begin
    int_issue_slot_5_com_1 = 12'h0;
    int_issue_slot_5_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_5.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_5.io_valid && !(soc1.core.int_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_5.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_5.slot_uop_rob_idx))
      begin
        int_issue_slot_5_com_1 = soc1.core.int_issue_unit.slots_5.slot_uop_br_mask;
        int_issue_slot_5_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_5_com_1 = 12'h0;
        int_issue_slot_5_uncom_1 = soc1.core.int_issue_unit.slots_5.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_6_com_1;
  wire [11:0] int_issue_slot_6_uncom_1;

  always @(*)
  begin
    int_issue_slot_6_com_1 = 12'h0;
    int_issue_slot_6_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_6.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_6.io_valid && !(soc1.core.int_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_6.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_6.slot_uop_rob_idx))
      begin
        int_issue_slot_6_com_1 = soc1.core.int_issue_unit.slots_6.slot_uop_br_mask;
        int_issue_slot_6_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_6_com_1 = 12'h0;
        int_issue_slot_6_uncom_1 = soc1.core.int_issue_unit.slots_6.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_7_com_1;
  wire [11:0] int_issue_slot_7_uncom_1;

  always @(*)
  begin
    int_issue_slot_7_com_1 = 12'h0;
    int_issue_slot_7_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_7.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_7.io_valid && !(soc1.core.int_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_7.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_7.slot_uop_rob_idx))
      begin
        int_issue_slot_7_com_1 = soc1.core.int_issue_unit.slots_7.slot_uop_br_mask;
        int_issue_slot_7_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_7_com_1 = 12'h0;
        int_issue_slot_7_uncom_1 = soc1.core.int_issue_unit.slots_7.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_8_com_1;
  wire [11:0] int_issue_slot_8_uncom_1;

  always @(*)
  begin
    int_issue_slot_8_com_1 = 12'h0;
    int_issue_slot_8_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_8.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_8.io_valid && !(soc1.core.int_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_8.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_8.slot_uop_rob_idx))
      begin
        int_issue_slot_8_com_1 = soc1.core.int_issue_unit.slots_8.slot_uop_br_mask;
        int_issue_slot_8_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_8_com_1 = 12'h0;
        int_issue_slot_8_uncom_1 = soc1.core.int_issue_unit.slots_8.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_9_com_1;
  wire [11:0] int_issue_slot_9_uncom_1;

  always @(*)
  begin
    int_issue_slot_9_com_1 = 12'h0;
    int_issue_slot_9_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_9.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_9.io_valid && !(soc1.core.int_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_9.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_9.slot_uop_rob_idx))
      begin
        int_issue_slot_9_com_1 = soc1.core.int_issue_unit.slots_9.slot_uop_br_mask;
        int_issue_slot_9_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_9_com_1 = 12'h0;
        int_issue_slot_9_uncom_1 = soc1.core.int_issue_unit.slots_9.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_10_com_1;
  wire [11:0] int_issue_slot_10_uncom_1;

  always @(*)
  begin
    int_issue_slot_10_com_1 = 12'h0;
    int_issue_slot_10_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_10.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_10.io_valid && !(soc1.core.int_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_10.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_10.slot_uop_rob_idx))
      begin
        int_issue_slot_10_com_1 = soc1.core.int_issue_unit.slots_10.slot_uop_br_mask;
        int_issue_slot_10_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_10_com_1 = 12'h0;
        int_issue_slot_10_uncom_1 = soc1.core.int_issue_unit.slots_10.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_11_com_1;
  wire [11:0] int_issue_slot_11_uncom_1;

  always @(*)
  begin
    int_issue_slot_11_com_1 = 12'h0;
    int_issue_slot_11_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_11.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_11.io_valid && !(soc1.core.int_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_11.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_11.slot_uop_rob_idx))
      begin
        int_issue_slot_11_com_1 = soc1.core.int_issue_unit.slots_11.slot_uop_br_mask;
        int_issue_slot_11_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_11_com_1 = 12'h0;
        int_issue_slot_11_uncom_1 = soc1.core.int_issue_unit.slots_11.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_12_com_1;
  wire [11:0] int_issue_slot_12_uncom_1;

  always @(*)
  begin
    int_issue_slot_12_com_1 = 12'h0;
    int_issue_slot_12_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_12.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_12.io_valid && !(soc1.core.int_issue_unit.slots_12.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_12.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_12.slot_uop_rob_idx))
      begin
        int_issue_slot_12_com_1 = soc1.core.int_issue_unit.slots_12.slot_uop_br_mask;
        int_issue_slot_12_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_12_com_1 = 12'h0;
        int_issue_slot_12_uncom_1 = soc1.core.int_issue_unit.slots_12.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_13_com_1;
  wire [11:0] int_issue_slot_13_uncom_1;

  always @(*)
  begin
    int_issue_slot_13_com_1 = 12'h0;
    int_issue_slot_13_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_13.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_13.io_valid && !(soc1.core.int_issue_unit.slots_13.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_13.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_13.slot_uop_rob_idx))
      begin
        int_issue_slot_13_com_1 = soc1.core.int_issue_unit.slots_13.slot_uop_br_mask;
        int_issue_slot_13_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_13_com_1 = 12'h0;
        int_issue_slot_13_uncom_1 = soc1.core.int_issue_unit.slots_13.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_14_com_1;
  wire [11:0] int_issue_slot_14_uncom_1;

  always @(*)
  begin
    int_issue_slot_14_com_1 = 12'h0;
    int_issue_slot_14_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_14.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_14.io_valid && !(soc1.core.int_issue_unit.slots_14.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_14.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_14.slot_uop_rob_idx))
      begin
        int_issue_slot_14_com_1 = soc1.core.int_issue_unit.slots_14.slot_uop_br_mask;
        int_issue_slot_14_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_14_com_1 = 12'h0;
        int_issue_slot_14_uncom_1 = soc1.core.int_issue_unit.slots_14.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_15_com_1;
  wire [11:0] int_issue_slot_15_uncom_1;

  always @(*)
  begin
    int_issue_slot_15_com_1 = 12'h0;
    int_issue_slot_15_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_15.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_15.io_valid && !(soc1.core.int_issue_unit.slots_15.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_15.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_15.slot_uop_rob_idx))
      begin
        int_issue_slot_15_com_1 = soc1.core.int_issue_unit.slots_15.slot_uop_br_mask;
        int_issue_slot_15_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_15_com_1 = 12'h0;
        int_issue_slot_15_uncom_1 = soc1.core.int_issue_unit.slots_15.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_16_com_1;
  wire [11:0] int_issue_slot_16_uncom_1;

  always @(*)
  begin
    int_issue_slot_16_com_1 = 12'h0;
    int_issue_slot_16_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_16.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_16.io_valid && !(soc1.core.int_issue_unit.slots_16.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_16.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_16.slot_uop_rob_idx))
      begin
        int_issue_slot_16_com_1 = soc1.core.int_issue_unit.slots_16.slot_uop_br_mask;
        int_issue_slot_16_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_16_com_1 = 12'h0;
        int_issue_slot_16_uncom_1 = soc1.core.int_issue_unit.slots_16.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_17_com_1;
  wire [11:0] int_issue_slot_17_uncom_1;

  always @(*)
  begin
    int_issue_slot_17_com_1 = 12'h0;
    int_issue_slot_17_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_17.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_17.io_valid && !(soc1.core.int_issue_unit.slots_17.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_17.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_17.slot_uop_rob_idx))
      begin
        int_issue_slot_17_com_1 = soc1.core.int_issue_unit.slots_17.slot_uop_br_mask;
        int_issue_slot_17_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_17_com_1 = 12'h0;
        int_issue_slot_17_uncom_1 = soc1.core.int_issue_unit.slots_17.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_18_com_1;
  wire [11:0] int_issue_slot_18_uncom_1;

  always @(*)
  begin
    int_issue_slot_18_com_1 = 12'h0;
    int_issue_slot_18_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_18.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_18.io_valid && !(soc1.core.int_issue_unit.slots_18.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_18.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_18.slot_uop_rob_idx))
      begin
        int_issue_slot_18_com_1 = soc1.core.int_issue_unit.slots_18.slot_uop_br_mask;
        int_issue_slot_18_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_18_com_1 = 12'h0;
        int_issue_slot_18_uncom_1 = soc1.core.int_issue_unit.slots_18.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_19_com_1;
  wire [11:0] int_issue_slot_19_uncom_1;

  always @(*)
  begin
    int_issue_slot_19_com_1 = 12'h0;
    int_issue_slot_19_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.int_issue_unit.slots_19.slot_uop_rob_idx) && soc1.core.int_issue_unit.slots_19.io_valid && !(soc1.core.int_issue_unit.slots_19.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_19.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_19.slot_uop_rob_idx))
      begin
        int_issue_slot_19_com_1 = soc1.core.int_issue_unit.slots_19.slot_uop_br_mask;
        int_issue_slot_19_uncom_1 = 12'hfff;
      end
      else
      begin
        int_issue_slot_19_com_1 = 12'h0;
        int_issue_slot_19_uncom_1 = soc1.core.int_issue_unit.slots_19.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_0_com_1;
  wire [11:0] mem_issue_slot_0_uncom_1;

  always @(*)
  begin
    mem_issue_slot_0_com_1 = 12'h0;
    mem_issue_slot_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_0.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_0.io_valid && !(soc1.core.mem_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_0.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_0.slot_uop_rob_idx))
      begin
        mem_issue_slot_0_com_1 = soc1.core.mem_issue_unit.slots_0.slot_uop_br_mask;
        mem_issue_slot_0_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_0_com_1 = 12'h0;
        mem_issue_slot_0_uncom_1 = soc1.core.mem_issue_unit.slots_0.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_1_com_1;
  wire [11:0] mem_issue_slot_1_uncom_1;

  always @(*)
  begin
    mem_issue_slot_1_com_1 = 12'h0;
    mem_issue_slot_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_1.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_1.io_valid && !(soc1.core.mem_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_1.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_1.slot_uop_rob_idx))
      begin
        mem_issue_slot_1_com_1 = soc1.core.mem_issue_unit.slots_1.slot_uop_br_mask;
        mem_issue_slot_1_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_1_com_1 = 12'h0;
        mem_issue_slot_1_uncom_1 = soc1.core.mem_issue_unit.slots_1.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_2_com_1;
  wire [11:0] mem_issue_slot_2_uncom_1;

  always @(*)
  begin
    mem_issue_slot_2_com_1 = 12'h0;
    mem_issue_slot_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_2.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_2.io_valid && !(soc1.core.mem_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_2.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_2.slot_uop_rob_idx))
      begin
        mem_issue_slot_2_com_1 = soc1.core.mem_issue_unit.slots_2.slot_uop_br_mask;
        mem_issue_slot_2_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_2_com_1 = 12'h0;
        mem_issue_slot_2_uncom_1 = soc1.core.mem_issue_unit.slots_2.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_3_com_1;
  wire [11:0] mem_issue_slot_3_uncom_1;

  always @(*)
  begin
    mem_issue_slot_3_com_1 = 12'h0;
    mem_issue_slot_3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_3.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_3.io_valid && !(soc1.core.mem_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_3.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_3.slot_uop_rob_idx))
      begin
        mem_issue_slot_3_com_1 = soc1.core.mem_issue_unit.slots_3.slot_uop_br_mask;
        mem_issue_slot_3_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_3_com_1 = 12'h0;
        mem_issue_slot_3_uncom_1 = soc1.core.mem_issue_unit.slots_3.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_4_com_1;
  wire [11:0] mem_issue_slot_4_uncom_1;

  always @(*)
  begin
    mem_issue_slot_4_com_1 = 12'h0;
    mem_issue_slot_4_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_4.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_4.io_valid && !(soc1.core.mem_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_4.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_4.slot_uop_rob_idx))
      begin
        mem_issue_slot_4_com_1 = soc1.core.mem_issue_unit.slots_4.slot_uop_br_mask;
        mem_issue_slot_4_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_4_com_1 = 12'h0;
        mem_issue_slot_4_uncom_1 = soc1.core.mem_issue_unit.slots_4.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_5_com_1;
  wire [11:0] mem_issue_slot_5_uncom_1;

  always @(*)
  begin
    mem_issue_slot_5_com_1 = 12'h0;
    mem_issue_slot_5_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_5.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_5.io_valid && !(soc1.core.mem_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_5.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_5.slot_uop_rob_idx))
      begin
        mem_issue_slot_5_com_1 = soc1.core.mem_issue_unit.slots_5.slot_uop_br_mask;
        mem_issue_slot_5_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_5_com_1 = 12'h0;
        mem_issue_slot_5_uncom_1 = soc1.core.mem_issue_unit.slots_5.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_6_com_1;
  wire [11:0] mem_issue_slot_6_uncom_1;

  always @(*)
  begin
    mem_issue_slot_6_com_1 = 12'h0;
    mem_issue_slot_6_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_6.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_6.io_valid && !(soc1.core.mem_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_6.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_6.slot_uop_rob_idx))
      begin
        mem_issue_slot_6_com_1 = soc1.core.mem_issue_unit.slots_6.slot_uop_br_mask;
        mem_issue_slot_6_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_6_com_1 = 12'h0;
        mem_issue_slot_6_uncom_1 = soc1.core.mem_issue_unit.slots_6.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_7_com_1;
  wire [11:0] mem_issue_slot_7_uncom_1;

  always @(*)
  begin
    mem_issue_slot_7_com_1 = 12'h0;
    mem_issue_slot_7_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_7.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_7.io_valid && !(soc1.core.mem_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_7.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_7.slot_uop_rob_idx))
      begin
        mem_issue_slot_7_com_1 = soc1.core.mem_issue_unit.slots_7.slot_uop_br_mask;
        mem_issue_slot_7_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_7_com_1 = 12'h0;
        mem_issue_slot_7_uncom_1 = soc1.core.mem_issue_unit.slots_7.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_8_com_1;
  wire [11:0] mem_issue_slot_8_uncom_1;

  always @(*)
  begin
    mem_issue_slot_8_com_1 = 12'h0;
    mem_issue_slot_8_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_8.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_8.io_valid && !(soc1.core.mem_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_8.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_8.slot_uop_rob_idx))
      begin
        mem_issue_slot_8_com_1 = soc1.core.mem_issue_unit.slots_8.slot_uop_br_mask;
        mem_issue_slot_8_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_8_com_1 = 12'h0;
        mem_issue_slot_8_uncom_1 = soc1.core.mem_issue_unit.slots_8.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_9_com_1;
  wire [11:0] mem_issue_slot_9_uncom_1;

  always @(*)
  begin
    mem_issue_slot_9_com_1 = 12'h0;
    mem_issue_slot_9_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_9.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_9.io_valid && !(soc1.core.mem_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_9.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_9.slot_uop_rob_idx))
      begin
        mem_issue_slot_9_com_1 = soc1.core.mem_issue_unit.slots_9.slot_uop_br_mask;
        mem_issue_slot_9_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_9_com_1 = 12'h0;
        mem_issue_slot_9_uncom_1 = soc1.core.mem_issue_unit.slots_9.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_10_com_1;
  wire [11:0] mem_issue_slot_10_uncom_1;

  always @(*)
  begin
    mem_issue_slot_10_com_1 = 12'h0;
    mem_issue_slot_10_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_10.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_10.io_valid && !(soc1.core.mem_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_10.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_10.slot_uop_rob_idx))
      begin
        mem_issue_slot_10_com_1 = soc1.core.mem_issue_unit.slots_10.slot_uop_br_mask;
        mem_issue_slot_10_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_10_com_1 = 12'h0;
        mem_issue_slot_10_uncom_1 = soc1.core.mem_issue_unit.slots_10.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_11_com_1;
  wire [11:0] mem_issue_slot_11_uncom_1;

  always @(*)
  begin
    mem_issue_slot_11_com_1 = 12'h0;
    mem_issue_slot_11_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.core.mem_issue_unit.slots_11.slot_uop_rob_idx) && soc1.core.mem_issue_unit.slots_11.io_valid && !(soc1.core.mem_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_11.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_11.slot_uop_rob_idx))
      begin
        mem_issue_slot_11_com_1 = soc1.core.mem_issue_unit.slots_11.slot_uop_br_mask;
        mem_issue_slot_11_uncom_1 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_11_com_1 = 12'h0;
        mem_issue_slot_11_uncom_1 = soc1.core.mem_issue_unit.slots_11.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_0_com_1;
  wire [11:0] lsu_ldq_0_uncom_1;

  always @(*)
  begin
    lsu_ldq_0_com_1 = 12'h0;
    lsu_ldq_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_0_bits_uop_rob_idx) && soc1.lsu.ldq_0_valid && !(soc1.lsu.ldq_0_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_0_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_0_bits_uop_rob_idx))
      begin
        lsu_ldq_0_com_1 = soc1.lsu.ldq_0_bits_uop_br_mask;
        lsu_ldq_0_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_0_com_1 = 12'h0;
        lsu_ldq_0_uncom_1 = soc1.lsu.ldq_0_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_1_com_1;
  wire [11:0] lsu_ldq_1_uncom_1;

  always @(*)
  begin
    lsu_ldq_1_com_1 = 12'h0;
    lsu_ldq_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_1_bits_uop_rob_idx) && soc1.lsu.ldq_1_valid && !(soc1.lsu.ldq_1_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_1_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_1_bits_uop_rob_idx))
      begin
        lsu_ldq_1_com_1 = soc1.lsu.ldq_1_bits_uop_br_mask;
        lsu_ldq_1_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_1_com_1 = 12'h0;
        lsu_ldq_1_uncom_1 = soc1.lsu.ldq_1_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_2_com_1;
  wire [11:0] lsu_ldq_2_uncom_1;

  always @(*)
  begin
    lsu_ldq_2_com_1 = 12'h0;
    lsu_ldq_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_2_bits_uop_rob_idx) && soc1.lsu.ldq_2_valid && !(soc1.lsu.ldq_2_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_2_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_2_bits_uop_rob_idx))
      begin
        lsu_ldq_2_com_1 = soc1.lsu.ldq_2_bits_uop_br_mask;
        lsu_ldq_2_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_2_com_1 = 12'h0;
        lsu_ldq_2_uncom_1 = soc1.lsu.ldq_2_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_3_com_1;
  wire [11:0] lsu_ldq_3_uncom_1;

  always @(*)
  begin
    lsu_ldq_3_com_1 = 12'h0;
    lsu_ldq_3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_3_bits_uop_rob_idx) && soc1.lsu.ldq_3_valid && !(soc1.lsu.ldq_3_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_3_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_3_bits_uop_rob_idx))
      begin
        lsu_ldq_3_com_1 = soc1.lsu.ldq_3_bits_uop_br_mask;
        lsu_ldq_3_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_3_com_1 = 12'h0;
        lsu_ldq_3_uncom_1 = soc1.lsu.ldq_3_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_4_com_1;
  wire [11:0] lsu_ldq_4_uncom_1;

  always @(*)
  begin
    lsu_ldq_4_com_1 = 12'h0;
    lsu_ldq_4_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_4_bits_uop_rob_idx) && soc1.lsu.ldq_4_valid && !(soc1.lsu.ldq_4_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_4_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_4_bits_uop_rob_idx))
      begin
        lsu_ldq_4_com_1 = soc1.lsu.ldq_4_bits_uop_br_mask;
        lsu_ldq_4_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_4_com_1 = 12'h0;
        lsu_ldq_4_uncom_1 = soc1.lsu.ldq_4_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_5_com_1;
  wire [11:0] lsu_ldq_5_uncom_1;

  always @(*)
  begin
    lsu_ldq_5_com_1 = 12'h0;
    lsu_ldq_5_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_5_bits_uop_rob_idx) && soc1.lsu.ldq_5_valid && !(soc1.lsu.ldq_5_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_5_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_5_bits_uop_rob_idx))
      begin
        lsu_ldq_5_com_1 = soc1.lsu.ldq_5_bits_uop_br_mask;
        lsu_ldq_5_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_5_com_1 = 12'h0;
        lsu_ldq_5_uncom_1 = soc1.lsu.ldq_5_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_6_com_1;
  wire [11:0] lsu_ldq_6_uncom_1;

  always @(*)
  begin
    lsu_ldq_6_com_1 = 12'h0;
    lsu_ldq_6_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_6_bits_uop_rob_idx) && soc1.lsu.ldq_6_valid && !(soc1.lsu.ldq_6_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_6_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_6_bits_uop_rob_idx))
      begin
        lsu_ldq_6_com_1 = soc1.lsu.ldq_6_bits_uop_br_mask;
        lsu_ldq_6_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_6_com_1 = 12'h0;
        lsu_ldq_6_uncom_1 = soc1.lsu.ldq_6_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_7_com_1;
  wire [11:0] lsu_ldq_7_uncom_1;

  always @(*)
  begin
    lsu_ldq_7_com_1 = 12'h0;
    lsu_ldq_7_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_7_bits_uop_rob_idx) && soc1.lsu.ldq_7_valid && !(soc1.lsu.ldq_7_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_7_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_7_bits_uop_rob_idx))
      begin
        lsu_ldq_7_com_1 = soc1.lsu.ldq_7_bits_uop_br_mask;
        lsu_ldq_7_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_7_com_1 = 12'h0;
        lsu_ldq_7_uncom_1 = soc1.lsu.ldq_7_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_8_com_1;
  wire [11:0] lsu_ldq_8_uncom_1;

  always @(*)
  begin
    lsu_ldq_8_com_1 = 12'h0;
    lsu_ldq_8_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_8_bits_uop_rob_idx) && soc1.lsu.ldq_8_valid && !(soc1.lsu.ldq_8_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_8_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_8_bits_uop_rob_idx))
      begin
        lsu_ldq_8_com_1 = soc1.lsu.ldq_8_bits_uop_br_mask;
        lsu_ldq_8_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_8_com_1 = 12'h0;
        lsu_ldq_8_uncom_1 = soc1.lsu.ldq_8_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_9_com_1;
  wire [11:0] lsu_ldq_9_uncom_1;

  always @(*)
  begin
    lsu_ldq_9_com_1 = 12'h0;
    lsu_ldq_9_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_9_bits_uop_rob_idx) && soc1.lsu.ldq_9_valid && !(soc1.lsu.ldq_9_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_9_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_9_bits_uop_rob_idx))
      begin
        lsu_ldq_9_com_1 = soc1.lsu.ldq_9_bits_uop_br_mask;
        lsu_ldq_9_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_9_com_1 = 12'h0;
        lsu_ldq_9_uncom_1 = soc1.lsu.ldq_9_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_10_com_1;
  wire [11:0] lsu_ldq_10_uncom_1;

  always @(*)
  begin
    lsu_ldq_10_com_1 = 12'h0;
    lsu_ldq_10_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_10_bits_uop_rob_idx) && soc1.lsu.ldq_10_valid && !(soc1.lsu.ldq_10_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_10_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_10_bits_uop_rob_idx))
      begin
        lsu_ldq_10_com_1 = soc1.lsu.ldq_10_bits_uop_br_mask;
        lsu_ldq_10_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_10_com_1 = 12'h0;
        lsu_ldq_10_uncom_1 = soc1.lsu.ldq_10_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_11_com_1;
  wire [11:0] lsu_ldq_11_uncom_1;

  always @(*)
  begin
    lsu_ldq_11_com_1 = 12'h0;
    lsu_ldq_11_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_11_bits_uop_rob_idx) && soc1.lsu.ldq_11_valid && !(soc1.lsu.ldq_11_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_11_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_11_bits_uop_rob_idx))
      begin
        lsu_ldq_11_com_1 = soc1.lsu.ldq_11_bits_uop_br_mask;
        lsu_ldq_11_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_11_com_1 = 12'h0;
        lsu_ldq_11_uncom_1 = soc1.lsu.ldq_11_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_12_com_1;
  wire [11:0] lsu_ldq_12_uncom_1;

  always @(*)
  begin
    lsu_ldq_12_com_1 = 12'h0;
    lsu_ldq_12_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_12_bits_uop_rob_idx) && soc1.lsu.ldq_12_valid && !(soc1.lsu.ldq_12_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_12_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_12_bits_uop_rob_idx))
      begin
        lsu_ldq_12_com_1 = soc1.lsu.ldq_12_bits_uop_br_mask;
        lsu_ldq_12_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_12_com_1 = 12'h0;
        lsu_ldq_12_uncom_1 = soc1.lsu.ldq_12_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_13_com_1;
  wire [11:0] lsu_ldq_13_uncom_1;

  always @(*)
  begin
    lsu_ldq_13_com_1 = 12'h0;
    lsu_ldq_13_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_13_bits_uop_rob_idx) && soc1.lsu.ldq_13_valid && !(soc1.lsu.ldq_13_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_13_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_13_bits_uop_rob_idx))
      begin
        lsu_ldq_13_com_1 = soc1.lsu.ldq_13_bits_uop_br_mask;
        lsu_ldq_13_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_13_com_1 = 12'h0;
        lsu_ldq_13_uncom_1 = soc1.lsu.ldq_13_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_14_com_1;
  wire [11:0] lsu_ldq_14_uncom_1;

  always @(*)
  begin
    lsu_ldq_14_com_1 = 12'h0;
    lsu_ldq_14_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_14_bits_uop_rob_idx) && soc1.lsu.ldq_14_valid && !(soc1.lsu.ldq_14_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_14_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_14_bits_uop_rob_idx))
      begin
        lsu_ldq_14_com_1 = soc1.lsu.ldq_14_bits_uop_br_mask;
        lsu_ldq_14_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_14_com_1 = 12'h0;
        lsu_ldq_14_uncom_1 = soc1.lsu.ldq_14_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_15_com_1;
  wire [11:0] lsu_ldq_15_uncom_1;

  always @(*)
  begin
    lsu_ldq_15_com_1 = 12'h0;
    lsu_ldq_15_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.ldq_15_bits_uop_rob_idx) && soc1.lsu.ldq_15_valid && !(soc1.lsu.ldq_15_bits_uop_uses_stq && stq_committed_1[soc1.lsu.ldq_15_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_15_bits_uop_rob_idx))
      begin
        lsu_ldq_15_com_1 = soc1.lsu.ldq_15_bits_uop_br_mask;
        lsu_ldq_15_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_ldq_15_com_1 = 12'h0;
        lsu_ldq_15_uncom_1 = soc1.lsu.ldq_15_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_com_1;
  wire [11:0] lsu_mem_uncom_1;

  always @(*)
  begin
    lsu_mem_com_1 = 12'h0;
    lsu_mem_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.mem_incoming_uop_0_rob_idx) && soc1.lsu.fired_sfence_0)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.mem_incoming_uop_0_rob_idx))
      begin
        lsu_mem_com_1 = soc1.lsu.mem_incoming_uop_0_br_mask;
        lsu_mem_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_mem_com_1 = 12'h0;
        lsu_mem_uncom_1 = soc1.lsu.mem_incoming_uop_0_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_stq_com_1;
  wire [11:0] lsu_mem_stq_uncom_1;

  always @(*)
  begin
    lsu_mem_stq_com_1 = 12'h0;
    lsu_mem_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx) && (soc1.lsu.fired_stad_incoming_REG || soc1.lsu.fired_sta_incoming_REG || soc1.lsu.fired_std_incoming_REG) && !(stq_committed_1[soc1.lsu.mem_stq_incoming_e_0_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx))
      begin
        lsu_mem_stq_com_1 = soc1.lsu.mem_stq_incoming_e_0_bits_uop_br_mask;
        lsu_mem_stq_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_mem_stq_com_1 = 12'h0;
        lsu_mem_stq_uncom_1 = soc1.lsu.mem_stq_incoming_e_0_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_retry_com_1;
  wire [11:0] lsu_mem_retry_uncom_1;

  always @(*)
  begin
    lsu_mem_retry_com_1 = 12'h0;
    lsu_mem_retry_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.mem_stq_retry_e_bits_uop_rob_idx) && soc1.lsu.fired_sta_retry_REG && !(stq_committed_1[soc1.lsu.mem_stq_retry_e_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.mem_stq_retry_e_bits_uop_rob_idx))
      begin
        lsu_mem_retry_com_1 = soc1.lsu.mem_stq_retry_e_bits_uop_br_mask;
        lsu_mem_retry_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_mem_retry_com_1 = 12'h0;
        lsu_mem_retry_uncom_1 = soc1.lsu.mem_stq_retry_e_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_xcpt_com_1;
  wire [11:0] lsu_mem_xcpt_uncom_1;

  always @(*)
  begin
    lsu_mem_xcpt_com_1 = 12'h0;
    lsu_mem_xcpt_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.mem_xcpt_uops_0_rob_idx) && soc1.lsu.mem_xcpt_valids_0 && !(soc1.lsu.mem_xcpt_uops_0_uses_stq && stq_committed_1[soc1.lsu.mem_xcpt_uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.mem_xcpt_uops_0_rob_idx))
      begin
        lsu_mem_xcpt_com_1 = soc1.lsu.mem_xcpt_uops_0_br_mask;
        lsu_mem_xcpt_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_mem_xcpt_com_1 = 12'h0;
        lsu_mem_xcpt_uncom_1 = soc1.lsu.mem_xcpt_uops_0_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_stdf_com_1;
  wire [11:0] lsu_mem_stdf_uncom_1;

  always @(*)
  begin
    lsu_mem_stdf_com_1 = 12'h0;
    lsu_mem_stdf_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.mem_stdf_uop_rob_idx) && soc1.lsu.fired_stdf_incoming && !(stq_committed_1[soc1.lsu.mem_stdf_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.mem_stdf_uop_rob_idx))
      begin
        lsu_mem_stdf_com_1 = soc1.lsu.mem_stdf_uop_br_mask;
        lsu_mem_stdf_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_mem_stdf_com_1 = 12'h0;
        lsu_mem_stdf_uncom_1 = soc1.lsu.mem_stdf_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stdf_com_1;
  wire [11:0] lsu_stdf_uncom_1;

  always @(*)
  begin
    lsu_stdf_com_1 = 12'h0;
    lsu_stdf_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stdf_clr_bsy_rob_idx) && soc1.lsu.stdf_clr_bsy_valid)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stdf_clr_bsy_rob_idx))
      begin
        lsu_stdf_com_1 = soc1.lsu.stdf_clr_bsy_brmask;
        lsu_stdf_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stdf_com_1 = 12'h0;
        lsu_stdf_uncom_1 = soc1.lsu.stdf_clr_bsy_brmask;
      end
    end
  end

  wire [11:0] lsu_stq_0_com_1;
  wire [11:0] lsu_stq_0_uncom_1;

  always @(*)
  begin
    lsu_stq_0_com_1 = 12'h0;
    lsu_stq_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_0_bits_uop_rob_idx) && soc1.lsu.stq_0_valid && !soc1.lsu.stq_0_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_0_bits_uop_rob_idx))
      begin
        lsu_stq_0_com_1 = soc1.lsu.stq_0_bits_uop_br_mask;
        lsu_stq_0_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_0_com_1 = 12'h0;
        lsu_stq_0_uncom_1 = soc1.lsu.stq_0_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_1_com_1;
  wire [11:0] lsu_stq_1_uncom_1;

  always @(*)
  begin
    lsu_stq_1_com_1 = 12'h0;
    lsu_stq_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_1_bits_uop_rob_idx) && soc1.lsu.stq_1_valid && !soc1.lsu.stq_1_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_1_bits_uop_rob_idx))
      begin
        lsu_stq_1_com_1 = soc1.lsu.stq_1_bits_uop_br_mask;
        lsu_stq_1_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_1_com_1 = 12'h0;
        lsu_stq_1_uncom_1 = soc1.lsu.stq_1_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_2_com_1;
  wire [11:0] lsu_stq_2_uncom_1;

  always @(*)
  begin
    lsu_stq_2_com_1 = 12'h0;
    lsu_stq_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_2_bits_uop_rob_idx) && soc1.lsu.stq_2_valid && !soc1.lsu.stq_2_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_2_bits_uop_rob_idx))
      begin
        lsu_stq_2_com_1 = soc1.lsu.stq_2_bits_uop_br_mask;
        lsu_stq_2_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_2_com_1 = 12'h0;
        lsu_stq_2_uncom_1 = soc1.lsu.stq_2_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_3_com_1;
  wire [11:0] lsu_stq_3_uncom_1;

  always @(*)
  begin
    lsu_stq_3_com_1 = 12'h0;
    lsu_stq_3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_3_bits_uop_rob_idx) && soc1.lsu.stq_3_valid && !soc1.lsu.stq_3_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_3_bits_uop_rob_idx))
      begin
        lsu_stq_3_com_1 = soc1.lsu.stq_3_bits_uop_br_mask;
        lsu_stq_3_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_3_com_1 = 12'h0;
        lsu_stq_3_uncom_1 = soc1.lsu.stq_3_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_4_com_1;
  wire [11:0] lsu_stq_4_uncom_1;

  always @(*)
  begin
    lsu_stq_4_com_1 = 12'h0;
    lsu_stq_4_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_4_bits_uop_rob_idx) && soc1.lsu.stq_4_valid && !soc1.lsu.stq_4_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_4_bits_uop_rob_idx))
      begin
        lsu_stq_4_com_1 = soc1.lsu.stq_4_bits_uop_br_mask;
        lsu_stq_4_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_4_com_1 = 12'h0;
        lsu_stq_4_uncom_1 = soc1.lsu.stq_4_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_5_com_1;
  wire [11:0] lsu_stq_5_uncom_1;

  always @(*)
  begin
    lsu_stq_5_com_1 = 12'h0;
    lsu_stq_5_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_5_bits_uop_rob_idx) && soc1.lsu.stq_5_valid && !soc1.lsu.stq_5_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_5_bits_uop_rob_idx))
      begin
        lsu_stq_5_com_1 = soc1.lsu.stq_5_bits_uop_br_mask;
        lsu_stq_5_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_5_com_1 = 12'h0;
        lsu_stq_5_uncom_1 = soc1.lsu.stq_5_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_6_com_1;
  wire [11:0] lsu_stq_6_uncom_1;

  always @(*)
  begin
    lsu_stq_6_com_1 = 12'h0;
    lsu_stq_6_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_6_bits_uop_rob_idx) && soc1.lsu.stq_6_valid && !soc1.lsu.stq_6_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_6_bits_uop_rob_idx))
      begin
        lsu_stq_6_com_1 = soc1.lsu.stq_6_bits_uop_br_mask;
        lsu_stq_6_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_6_com_1 = 12'h0;
        lsu_stq_6_uncom_1 = soc1.lsu.stq_6_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_7_com_1;
  wire [11:0] lsu_stq_7_uncom_1;

  always @(*)
  begin
    lsu_stq_7_com_1 = 12'h0;
    lsu_stq_7_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_7_bits_uop_rob_idx) && soc1.lsu.stq_7_valid && !soc1.lsu.stq_7_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_7_bits_uop_rob_idx))
      begin
        lsu_stq_7_com_1 = soc1.lsu.stq_7_bits_uop_br_mask;
        lsu_stq_7_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_7_com_1 = 12'h0;
        lsu_stq_7_uncom_1 = soc1.lsu.stq_7_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_8_com_1;
  wire [11:0] lsu_stq_8_uncom_1;

  always @(*)
  begin
    lsu_stq_8_com_1 = 12'h0;
    lsu_stq_8_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_8_bits_uop_rob_idx) && soc1.lsu.stq_8_valid && !soc1.lsu.stq_8_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_8_bits_uop_rob_idx))
      begin
        lsu_stq_8_com_1 = soc1.lsu.stq_8_bits_uop_br_mask;
        lsu_stq_8_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_8_com_1 = 12'h0;
        lsu_stq_8_uncom_1 = soc1.lsu.stq_8_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_9_com_1;
  wire [11:0] lsu_stq_9_uncom_1;

  always @(*)
  begin
    lsu_stq_9_com_1 = 12'h0;
    lsu_stq_9_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_9_bits_uop_rob_idx) && soc1.lsu.stq_9_valid && !soc1.lsu.stq_9_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_9_bits_uop_rob_idx))
      begin
        lsu_stq_9_com_1 = soc1.lsu.stq_9_bits_uop_br_mask;
        lsu_stq_9_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_9_com_1 = 12'h0;
        lsu_stq_9_uncom_1 = soc1.lsu.stq_9_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_10_com_1;
  wire [11:0] lsu_stq_10_uncom_1;

  always @(*)
  begin
    lsu_stq_10_com_1 = 12'h0;
    lsu_stq_10_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_10_bits_uop_rob_idx) && soc1.lsu.stq_10_valid && !soc1.lsu.stq_10_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_10_bits_uop_rob_idx))
      begin
        lsu_stq_10_com_1 = soc1.lsu.stq_10_bits_uop_br_mask;
        lsu_stq_10_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_10_com_1 = 12'h0;
        lsu_stq_10_uncom_1 = soc1.lsu.stq_10_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_11_com_1;
  wire [11:0] lsu_stq_11_uncom_1;

  always @(*)
  begin
    lsu_stq_11_com_1 = 12'h0;
    lsu_stq_11_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_11_bits_uop_rob_idx) && soc1.lsu.stq_11_valid && !soc1.lsu.stq_11_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_11_bits_uop_rob_idx))
      begin
        lsu_stq_11_com_1 = soc1.lsu.stq_11_bits_uop_br_mask;
        lsu_stq_11_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_11_com_1 = 12'h0;
        lsu_stq_11_uncom_1 = soc1.lsu.stq_11_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_12_com_1;
  wire [11:0] lsu_stq_12_uncom_1;

  always @(*)
  begin
    lsu_stq_12_com_1 = 12'h0;
    lsu_stq_12_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_12_bits_uop_rob_idx) && soc1.lsu.stq_12_valid && !soc1.lsu.stq_12_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_12_bits_uop_rob_idx))
      begin
        lsu_stq_12_com_1 = soc1.lsu.stq_12_bits_uop_br_mask;
        lsu_stq_12_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_12_com_1 = 12'h0;
        lsu_stq_12_uncom_1 = soc1.lsu.stq_12_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_13_com_1;
  wire [11:0] lsu_stq_13_uncom_1;

  always @(*)
  begin
    lsu_stq_13_com_1 = 12'h0;
    lsu_stq_13_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_13_bits_uop_rob_idx) && soc1.lsu.stq_13_valid && !soc1.lsu.stq_13_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_13_bits_uop_rob_idx))
      begin
        lsu_stq_13_com_1 = soc1.lsu.stq_13_bits_uop_br_mask;
        lsu_stq_13_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_13_com_1 = 12'h0;
        lsu_stq_13_uncom_1 = soc1.lsu.stq_13_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_14_com_1;
  wire [11:0] lsu_stq_14_uncom_1;

  always @(*)
  begin
    lsu_stq_14_com_1 = 12'h0;
    lsu_stq_14_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_14_bits_uop_rob_idx) && soc1.lsu.stq_14_valid && !soc1.lsu.stq_14_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_14_bits_uop_rob_idx))
      begin
        lsu_stq_14_com_1 = soc1.lsu.stq_14_bits_uop_br_mask;
        lsu_stq_14_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_14_com_1 = 12'h0;
        lsu_stq_14_uncom_1 = soc1.lsu.stq_14_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_15_com_1;
  wire [11:0] lsu_stq_15_uncom_1;

  always @(*)
  begin
    lsu_stq_15_com_1 = 12'h0;
    lsu_stq_15_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.stq_15_bits_uop_rob_idx) && soc1.lsu.stq_15_valid && !soc1.lsu.stq_15_bits_committed)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_15_bits_uop_rob_idx))
      begin
        lsu_stq_15_com_1 = soc1.lsu.stq_15_bits_uop_br_mask;
        lsu_stq_15_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_stq_15_com_1 = 12'h0;
        lsu_stq_15_uncom_1 = soc1.lsu.stq_15_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] rob__0_com_1;
  wire [11:0] rob__0_uncom_1;

  always @(*)
  begin
    rob__0_com_1 = 12'h0;
    rob__0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b000000))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000000))
      begin
        rob__0_com_1 = soc1.core.rob.rob_uop__0_br_mask;
        rob__0_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__0_com_1 = 12'h0;
        rob__0_uncom_1 = soc1.core.rob.rob_uop__0_br_mask;
      end
    end
  end

  wire [11:0] rob__1_com_1;
  wire [11:0] rob__1_uncom_1;

  always @(*)
  begin
    rob__1_com_1 = 12'h0;
    rob__1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b000010))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000010))
      begin
        rob__1_com_1 = soc1.core.rob.rob_uop__1_br_mask;
        rob__1_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__1_com_1 = 12'h0;
        rob__1_uncom_1 = soc1.core.rob.rob_uop__1_br_mask;
      end
    end
  end

  wire [11:0] rob__2_com_1;
  wire [11:0] rob__2_uncom_1;

  always @(*)
  begin
    rob__2_com_1 = 12'h0;
    rob__2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b000100))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000100))
      begin
        rob__2_com_1 = soc1.core.rob.rob_uop__2_br_mask;
        rob__2_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__2_com_1 = 12'h0;
        rob__2_uncom_1 = soc1.core.rob.rob_uop__2_br_mask;
      end
    end
  end

  wire [11:0] rob__3_com_1;
  wire [11:0] rob__3_uncom_1;

  always @(*)
  begin
    rob__3_com_1 = 12'h0;
    rob__3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b000110))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000110))
      begin
        rob__3_com_1 = soc1.core.rob.rob_uop__3_br_mask;
        rob__3_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__3_com_1 = 12'h0;
        rob__3_uncom_1 = soc1.core.rob.rob_uop__3_br_mask;
      end
    end
  end

  wire [11:0] rob__4_com_1;
  wire [11:0] rob__4_uncom_1;

  always @(*)
  begin
    rob__4_com_1 = 12'h0;
    rob__4_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b001000))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001000))
      begin
        rob__4_com_1 = soc1.core.rob.rob_uop__4_br_mask;
        rob__4_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__4_com_1 = 12'h0;
        rob__4_uncom_1 = soc1.core.rob.rob_uop__4_br_mask;
      end
    end
  end

  wire [11:0] rob__5_com_1;
  wire [11:0] rob__5_uncom_1;

  always @(*)
  begin
    rob__5_com_1 = 12'h0;
    rob__5_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b001010))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001010))
      begin
        rob__5_com_1 = soc1.core.rob.rob_uop__5_br_mask;
        rob__5_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__5_com_1 = 12'h0;
        rob__5_uncom_1 = soc1.core.rob.rob_uop__5_br_mask;
      end
    end
  end

  wire [11:0] rob__6_com_1;
  wire [11:0] rob__6_uncom_1;

  always @(*)
  begin
    rob__6_com_1 = 12'h0;
    rob__6_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b001100))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001100))
      begin
        rob__6_com_1 = soc1.core.rob.rob_uop__6_br_mask;
        rob__6_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__6_com_1 = 12'h0;
        rob__6_uncom_1 = soc1.core.rob.rob_uop__6_br_mask;
      end
    end
  end

  wire [11:0] rob__7_com_1;
  wire [11:0] rob__7_uncom_1;

  always @(*)
  begin
    rob__7_com_1 = 12'h0;
    rob__7_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b001110))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001110))
      begin
        rob__7_com_1 = soc1.core.rob.rob_uop__7_br_mask;
        rob__7_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__7_com_1 = 12'h0;
        rob__7_uncom_1 = soc1.core.rob.rob_uop__7_br_mask;
      end
    end
  end

  wire [11:0] rob__8_com_1;
  wire [11:0] rob__8_uncom_1;

  always @(*)
  begin
    rob__8_com_1 = 12'h0;
    rob__8_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b010000))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010000))
      begin
        rob__8_com_1 = soc1.core.rob.rob_uop__8_br_mask;
        rob__8_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__8_com_1 = 12'h0;
        rob__8_uncom_1 = soc1.core.rob.rob_uop__8_br_mask;
      end
    end
  end

  wire [11:0] rob__9_com_1;
  wire [11:0] rob__9_uncom_1;

  always @(*)
  begin
    rob__9_com_1 = 12'h0;
    rob__9_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b010010))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010010))
      begin
        rob__9_com_1 = soc1.core.rob.rob_uop__9_br_mask;
        rob__9_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__9_com_1 = 12'h0;
        rob__9_uncom_1 = soc1.core.rob.rob_uop__9_br_mask;
      end
    end
  end

  wire [11:0] rob__10_com_1;
  wire [11:0] rob__10_uncom_1;

  always @(*)
  begin
    rob__10_com_1 = 12'h0;
    rob__10_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b010100))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010100))
      begin
        rob__10_com_1 = soc1.core.rob.rob_uop__10_br_mask;
        rob__10_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__10_com_1 = 12'h0;
        rob__10_uncom_1 = soc1.core.rob.rob_uop__10_br_mask;
      end
    end
  end

  wire [11:0] rob__11_com_1;
  wire [11:0] rob__11_uncom_1;

  always @(*)
  begin
    rob__11_com_1 = 12'h0;
    rob__11_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b010110))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010110))
      begin
        rob__11_com_1 = soc1.core.rob.rob_uop__11_br_mask;
        rob__11_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__11_com_1 = 12'h0;
        rob__11_uncom_1 = soc1.core.rob.rob_uop__11_br_mask;
      end
    end
  end

  wire [11:0] rob__12_com_1;
  wire [11:0] rob__12_uncom_1;

  always @(*)
  begin
    rob__12_com_1 = 12'h0;
    rob__12_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b011000))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011000))
      begin
        rob__12_com_1 = soc1.core.rob.rob_uop__12_br_mask;
        rob__12_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__12_com_1 = 12'h0;
        rob__12_uncom_1 = soc1.core.rob.rob_uop__12_br_mask;
      end
    end
  end

  wire [11:0] rob__13_com_1;
  wire [11:0] rob__13_uncom_1;

  always @(*)
  begin
    rob__13_com_1 = 12'h0;
    rob__13_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b011010))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011010))
      begin
        rob__13_com_1 = soc1.core.rob.rob_uop__13_br_mask;
        rob__13_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__13_com_1 = 12'h0;
        rob__13_uncom_1 = soc1.core.rob.rob_uop__13_br_mask;
      end
    end
  end

  wire [11:0] rob__14_com_1;
  wire [11:0] rob__14_uncom_1;

  always @(*)
  begin
    rob__14_com_1 = 12'h0;
    rob__14_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b011100))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011100))
      begin
        rob__14_com_1 = soc1.core.rob.rob_uop__14_br_mask;
        rob__14_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__14_com_1 = 12'h0;
        rob__14_uncom_1 = soc1.core.rob.rob_uop__14_br_mask;
      end
    end
  end

  wire [11:0] rob__15_com_1;
  wire [11:0] rob__15_uncom_1;

  always @(*)
  begin
    rob__15_com_1 = 12'h0;
    rob__15_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b011110))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011110))
      begin
        rob__15_com_1 = soc1.core.rob.rob_uop__15_br_mask;
        rob__15_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__15_com_1 = 12'h0;
        rob__15_uncom_1 = soc1.core.rob.rob_uop__15_br_mask;
      end
    end
  end

  wire [11:0] rob__16_com_1;
  wire [11:0] rob__16_uncom_1;

  always @(*)
  begin
    rob__16_com_1 = 12'h0;
    rob__16_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b100000))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100000))
      begin
        rob__16_com_1 = soc1.core.rob.rob_uop__16_br_mask;
        rob__16_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__16_com_1 = 12'h0;
        rob__16_uncom_1 = soc1.core.rob.rob_uop__16_br_mask;
      end
    end
  end

  wire [11:0] rob__17_com_1;
  wire [11:0] rob__17_uncom_1;

  always @(*)
  begin
    rob__17_com_1 = 12'h0;
    rob__17_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b100010))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100010))
      begin
        rob__17_com_1 = soc1.core.rob.rob_uop__17_br_mask;
        rob__17_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__17_com_1 = 12'h0;
        rob__17_uncom_1 = soc1.core.rob.rob_uop__17_br_mask;
      end
    end
  end

  wire [11:0] rob__18_com_1;
  wire [11:0] rob__18_uncom_1;

  always @(*)
  begin
    rob__18_com_1 = 12'h0;
    rob__18_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b100100))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100100))
      begin
        rob__18_com_1 = soc1.core.rob.rob_uop__18_br_mask;
        rob__18_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__18_com_1 = 12'h0;
        rob__18_uncom_1 = soc1.core.rob.rob_uop__18_br_mask;
      end
    end
  end

  wire [11:0] rob__19_com_1;
  wire [11:0] rob__19_uncom_1;

  always @(*)
  begin
    rob__19_com_1 = 12'h0;
    rob__19_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b100110))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100110))
      begin
        rob__19_com_1 = soc1.core.rob.rob_uop__19_br_mask;
        rob__19_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__19_com_1 = 12'h0;
        rob__19_uncom_1 = soc1.core.rob.rob_uop__19_br_mask;
      end
    end
  end

  wire [11:0] rob__20_com_1;
  wire [11:0] rob__20_uncom_1;

  always @(*)
  begin
    rob__20_com_1 = 12'h0;
    rob__20_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b101000))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101000))
      begin
        rob__20_com_1 = soc1.core.rob.rob_uop__20_br_mask;
        rob__20_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__20_com_1 = 12'h0;
        rob__20_uncom_1 = soc1.core.rob.rob_uop__20_br_mask;
      end
    end
  end

  wire [11:0] rob__21_com_1;
  wire [11:0] rob__21_uncom_1;

  always @(*)
  begin
    rob__21_com_1 = 12'h0;
    rob__21_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b101010))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101010))
      begin
        rob__21_com_1 = soc1.core.rob.rob_uop__21_br_mask;
        rob__21_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__21_com_1 = 12'h0;
        rob__21_uncom_1 = soc1.core.rob.rob_uop__21_br_mask;
      end
    end
  end

  wire [11:0] rob__22_com_1;
  wire [11:0] rob__22_uncom_1;

  always @(*)
  begin
    rob__22_com_1 = 12'h0;
    rob__22_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b101100))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101100))
      begin
        rob__22_com_1 = soc1.core.rob.rob_uop__22_br_mask;
        rob__22_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__22_com_1 = 12'h0;
        rob__22_uncom_1 = soc1.core.rob.rob_uop__22_br_mask;
      end
    end
  end

  wire [11:0] rob__23_com_1;
  wire [11:0] rob__23_uncom_1;

  always @(*)
  begin
    rob__23_com_1 = 12'h0;
    rob__23_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b101110))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101110))
      begin
        rob__23_com_1 = soc1.core.rob.rob_uop__23_br_mask;
        rob__23_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__23_com_1 = 12'h0;
        rob__23_uncom_1 = soc1.core.rob.rob_uop__23_br_mask;
      end
    end
  end

  wire [11:0] rob__24_com_1;
  wire [11:0] rob__24_uncom_1;

  always @(*)
  begin
    rob__24_com_1 = 12'h0;
    rob__24_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b110000))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110000))
      begin
        rob__24_com_1 = soc1.core.rob.rob_uop__24_br_mask;
        rob__24_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__24_com_1 = 12'h0;
        rob__24_uncom_1 = soc1.core.rob.rob_uop__24_br_mask;
      end
    end
  end

  wire [11:0] rob__25_com_1;
  wire [11:0] rob__25_uncom_1;

  always @(*)
  begin
    rob__25_com_1 = 12'h0;
    rob__25_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b110010))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110010))
      begin
        rob__25_com_1 = soc1.core.rob.rob_uop__25_br_mask;
        rob__25_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__25_com_1 = 12'h0;
        rob__25_uncom_1 = soc1.core.rob.rob_uop__25_br_mask;
      end
    end
  end

  wire [11:0] rob__26_com_1;
  wire [11:0] rob__26_uncom_1;

  always @(*)
  begin
    rob__26_com_1 = 12'h0;
    rob__26_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b110100))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110100))
      begin
        rob__26_com_1 = soc1.core.rob.rob_uop__26_br_mask;
        rob__26_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__26_com_1 = 12'h0;
        rob__26_uncom_1 = soc1.core.rob.rob_uop__26_br_mask;
      end
    end
  end

  wire [11:0] rob__27_com_1;
  wire [11:0] rob__27_uncom_1;

  always @(*)
  begin
    rob__27_com_1 = 12'h0;
    rob__27_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b110110))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110110))
      begin
        rob__27_com_1 = soc1.core.rob.rob_uop__27_br_mask;
        rob__27_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__27_com_1 = 12'h0;
        rob__27_uncom_1 = soc1.core.rob.rob_uop__27_br_mask;
      end
    end
  end

  wire [11:0] rob__28_com_1;
  wire [11:0] rob__28_uncom_1;

  always @(*)
  begin
    rob__28_com_1 = 12'h0;
    rob__28_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b111000))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111000))
      begin
        rob__28_com_1 = soc1.core.rob.rob_uop__28_br_mask;
        rob__28_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__28_com_1 = 12'h0;
        rob__28_uncom_1 = soc1.core.rob.rob_uop__28_br_mask;
      end
    end
  end

  wire [11:0] rob__29_com_1;
  wire [11:0] rob__29_uncom_1;

  always @(*)
  begin
    rob__29_com_1 = 12'h0;
    rob__29_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b111010))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111010))
      begin
        rob__29_com_1 = soc1.core.rob.rob_uop__29_br_mask;
        rob__29_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__29_com_1 = 12'h0;
        rob__29_uncom_1 = soc1.core.rob.rob_uop__29_br_mask;
      end
    end
  end

  wire [11:0] rob__30_com_1;
  wire [11:0] rob__30_uncom_1;

  always @(*)
  begin
    rob__30_com_1 = 12'h0;
    rob__30_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b111100))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111100))
      begin
        rob__30_com_1 = soc1.core.rob.rob_uop__30_br_mask;
        rob__30_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__30_com_1 = 12'h0;
        rob__30_uncom_1 = soc1.core.rob.rob_uop__30_br_mask;
      end
    end
  end

  wire [11:0] rob__31_com_1;
  wire [11:0] rob__31_uncom_1;

  always @(*)
  begin
    rob__31_com_1 = 12'h0;
    rob__31_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b111110))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111110))
      begin
        rob__31_com_1 = soc1.core.rob.rob_uop__31_br_mask;
        rob__31_uncom_1 = 12'hfff;
      end
      else
      begin
        rob__31_com_1 = 12'h0;
        rob__31_uncom_1 = soc1.core.rob.rob_uop__31_br_mask;
      end
    end
  end

  wire [11:0] rob_1_0_com_1;
  wire [11:0] rob_1_0_uncom_1;

  always @(*)
  begin
    rob_1_0_com_1 = 12'h0;
    rob_1_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b000001))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000001))
      begin
        rob_1_0_com_1 = soc1.core.rob.rob_uop_1_0_br_mask;
        rob_1_0_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_0_com_1 = 12'h0;
        rob_1_0_uncom_1 = soc1.core.rob.rob_uop_1_0_br_mask;
      end
    end
  end

  wire [11:0] rob_1_1_com_1;
  wire [11:0] rob_1_1_uncom_1;

  always @(*)
  begin
    rob_1_1_com_1 = 12'h0;
    rob_1_1_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b000011))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000011))
      begin
        rob_1_1_com_1 = soc1.core.rob.rob_uop_1_1_br_mask;
        rob_1_1_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_1_com_1 = 12'h0;
        rob_1_1_uncom_1 = soc1.core.rob.rob_uop_1_1_br_mask;
      end
    end
  end

  wire [11:0] rob_1_2_com_1;
  wire [11:0] rob_1_2_uncom_1;

  always @(*)
  begin
    rob_1_2_com_1 = 12'h0;
    rob_1_2_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b000101))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000101))
      begin
        rob_1_2_com_1 = soc1.core.rob.rob_uop_1_2_br_mask;
        rob_1_2_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_2_com_1 = 12'h0;
        rob_1_2_uncom_1 = soc1.core.rob.rob_uop_1_2_br_mask;
      end
    end
  end

  wire [11:0] rob_1_3_com_1;
  wire [11:0] rob_1_3_uncom_1;

  always @(*)
  begin
    rob_1_3_com_1 = 12'h0;
    rob_1_3_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b000111))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b000111))
      begin
        rob_1_3_com_1 = soc1.core.rob.rob_uop_1_3_br_mask;
        rob_1_3_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_3_com_1 = 12'h0;
        rob_1_3_uncom_1 = soc1.core.rob.rob_uop_1_3_br_mask;
      end
    end
  end

  wire [11:0] rob_1_4_com_1;
  wire [11:0] rob_1_4_uncom_1;

  always @(*)
  begin
    rob_1_4_com_1 = 12'h0;
    rob_1_4_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b001001))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001001))
      begin
        rob_1_4_com_1 = soc1.core.rob.rob_uop_1_4_br_mask;
        rob_1_4_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_4_com_1 = 12'h0;
        rob_1_4_uncom_1 = soc1.core.rob.rob_uop_1_4_br_mask;
      end
    end
  end

  wire [11:0] rob_1_5_com_1;
  wire [11:0] rob_1_5_uncom_1;

  always @(*)
  begin
    rob_1_5_com_1 = 12'h0;
    rob_1_5_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b001011))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001011))
      begin
        rob_1_5_com_1 = soc1.core.rob.rob_uop_1_5_br_mask;
        rob_1_5_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_5_com_1 = 12'h0;
        rob_1_5_uncom_1 = soc1.core.rob.rob_uop_1_5_br_mask;
      end
    end
  end

  wire [11:0] rob_1_6_com_1;
  wire [11:0] rob_1_6_uncom_1;

  always @(*)
  begin
    rob_1_6_com_1 = 12'h0;
    rob_1_6_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b001101))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001101))
      begin
        rob_1_6_com_1 = soc1.core.rob.rob_uop_1_6_br_mask;
        rob_1_6_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_6_com_1 = 12'h0;
        rob_1_6_uncom_1 = soc1.core.rob.rob_uop_1_6_br_mask;
      end
    end
  end

  wire [11:0] rob_1_7_com_1;
  wire [11:0] rob_1_7_uncom_1;

  always @(*)
  begin
    rob_1_7_com_1 = 12'h0;
    rob_1_7_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b001111))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b001111))
      begin
        rob_1_7_com_1 = soc1.core.rob.rob_uop_1_7_br_mask;
        rob_1_7_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_7_com_1 = 12'h0;
        rob_1_7_uncom_1 = soc1.core.rob.rob_uop_1_7_br_mask;
      end
    end
  end

  wire [11:0] rob_1_8_com_1;
  wire [11:0] rob_1_8_uncom_1;

  always @(*)
  begin
    rob_1_8_com_1 = 12'h0;
    rob_1_8_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b010001))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010001))
      begin
        rob_1_8_com_1 = soc1.core.rob.rob_uop_1_8_br_mask;
        rob_1_8_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_8_com_1 = 12'h0;
        rob_1_8_uncom_1 = soc1.core.rob.rob_uop_1_8_br_mask;
      end
    end
  end

  wire [11:0] rob_1_9_com_1;
  wire [11:0] rob_1_9_uncom_1;

  always @(*)
  begin
    rob_1_9_com_1 = 12'h0;
    rob_1_9_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b010011))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010011))
      begin
        rob_1_9_com_1 = soc1.core.rob.rob_uop_1_9_br_mask;
        rob_1_9_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_9_com_1 = 12'h0;
        rob_1_9_uncom_1 = soc1.core.rob.rob_uop_1_9_br_mask;
      end
    end
  end

  wire [11:0] rob_1_10_com_1;
  wire [11:0] rob_1_10_uncom_1;

  always @(*)
  begin
    rob_1_10_com_1 = 12'h0;
    rob_1_10_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b010101))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010101))
      begin
        rob_1_10_com_1 = soc1.core.rob.rob_uop_1_10_br_mask;
        rob_1_10_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_10_com_1 = 12'h0;
        rob_1_10_uncom_1 = soc1.core.rob.rob_uop_1_10_br_mask;
      end
    end
  end

  wire [11:0] rob_1_11_com_1;
  wire [11:0] rob_1_11_uncom_1;

  always @(*)
  begin
    rob_1_11_com_1 = 12'h0;
    rob_1_11_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b010111))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b010111))
      begin
        rob_1_11_com_1 = soc1.core.rob.rob_uop_1_11_br_mask;
        rob_1_11_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_11_com_1 = 12'h0;
        rob_1_11_uncom_1 = soc1.core.rob.rob_uop_1_11_br_mask;
      end
    end
  end

  wire [11:0] rob_1_12_com_1;
  wire [11:0] rob_1_12_uncom_1;

  always @(*)
  begin
    rob_1_12_com_1 = 12'h0;
    rob_1_12_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b011001))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011001))
      begin
        rob_1_12_com_1 = soc1.core.rob.rob_uop_1_12_br_mask;
        rob_1_12_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_12_com_1 = 12'h0;
        rob_1_12_uncom_1 = soc1.core.rob.rob_uop_1_12_br_mask;
      end
    end
  end

  wire [11:0] rob_1_13_com_1;
  wire [11:0] rob_1_13_uncom_1;

  always @(*)
  begin
    rob_1_13_com_1 = 12'h0;
    rob_1_13_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b011011))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011011))
      begin
        rob_1_13_com_1 = soc1.core.rob.rob_uop_1_13_br_mask;
        rob_1_13_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_13_com_1 = 12'h0;
        rob_1_13_uncom_1 = soc1.core.rob.rob_uop_1_13_br_mask;
      end
    end
  end

  wire [11:0] rob_1_14_com_1;
  wire [11:0] rob_1_14_uncom_1;

  always @(*)
  begin
    rob_1_14_com_1 = 12'h0;
    rob_1_14_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b011101))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011101))
      begin
        rob_1_14_com_1 = soc1.core.rob.rob_uop_1_14_br_mask;
        rob_1_14_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_14_com_1 = 12'h0;
        rob_1_14_uncom_1 = soc1.core.rob.rob_uop_1_14_br_mask;
      end
    end
  end

  wire [11:0] rob_1_15_com_1;
  wire [11:0] rob_1_15_uncom_1;

  always @(*)
  begin
    rob_1_15_com_1 = 12'h0;
    rob_1_15_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b011111))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b011111))
      begin
        rob_1_15_com_1 = soc1.core.rob.rob_uop_1_15_br_mask;
        rob_1_15_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_15_com_1 = 12'h0;
        rob_1_15_uncom_1 = soc1.core.rob.rob_uop_1_15_br_mask;
      end
    end
  end

  wire [11:0] rob_1_16_com_1;
  wire [11:0] rob_1_16_uncom_1;

  always @(*)
  begin
    rob_1_16_com_1 = 12'h0;
    rob_1_16_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b100001))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100001))
      begin
        rob_1_16_com_1 = soc1.core.rob.rob_uop_1_16_br_mask;
        rob_1_16_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_16_com_1 = 12'h0;
        rob_1_16_uncom_1 = soc1.core.rob.rob_uop_1_16_br_mask;
      end
    end
  end

  wire [11:0] rob_1_17_com_1;
  wire [11:0] rob_1_17_uncom_1;

  always @(*)
  begin
    rob_1_17_com_1 = 12'h0;
    rob_1_17_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b100011))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100011))
      begin
        rob_1_17_com_1 = soc1.core.rob.rob_uop_1_17_br_mask;
        rob_1_17_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_17_com_1 = 12'h0;
        rob_1_17_uncom_1 = soc1.core.rob.rob_uop_1_17_br_mask;
      end
    end
  end

  wire [11:0] rob_1_18_com_1;
  wire [11:0] rob_1_18_uncom_1;

  always @(*)
  begin
    rob_1_18_com_1 = 12'h0;
    rob_1_18_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b100101))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100101))
      begin
        rob_1_18_com_1 = soc1.core.rob.rob_uop_1_18_br_mask;
        rob_1_18_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_18_com_1 = 12'h0;
        rob_1_18_uncom_1 = soc1.core.rob.rob_uop_1_18_br_mask;
      end
    end
  end

  wire [11:0] rob_1_19_com_1;
  wire [11:0] rob_1_19_uncom_1;

  always @(*)
  begin
    rob_1_19_com_1 = 12'h0;
    rob_1_19_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b100111))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b100111))
      begin
        rob_1_19_com_1 = soc1.core.rob.rob_uop_1_19_br_mask;
        rob_1_19_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_19_com_1 = 12'h0;
        rob_1_19_uncom_1 = soc1.core.rob.rob_uop_1_19_br_mask;
      end
    end
  end

  wire [11:0] rob_1_20_com_1;
  wire [11:0] rob_1_20_uncom_1;

  always @(*)
  begin
    rob_1_20_com_1 = 12'h0;
    rob_1_20_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b101001))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101001))
      begin
        rob_1_20_com_1 = soc1.core.rob.rob_uop_1_20_br_mask;
        rob_1_20_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_20_com_1 = 12'h0;
        rob_1_20_uncom_1 = soc1.core.rob.rob_uop_1_20_br_mask;
      end
    end
  end

  wire [11:0] rob_1_21_com_1;
  wire [11:0] rob_1_21_uncom_1;

  always @(*)
  begin
    rob_1_21_com_1 = 12'h0;
    rob_1_21_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b101011))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101011))
      begin
        rob_1_21_com_1 = soc1.core.rob.rob_uop_1_21_br_mask;
        rob_1_21_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_21_com_1 = 12'h0;
        rob_1_21_uncom_1 = soc1.core.rob.rob_uop_1_21_br_mask;
      end
    end
  end

  wire [11:0] rob_1_22_com_1;
  wire [11:0] rob_1_22_uncom_1;

  always @(*)
  begin
    rob_1_22_com_1 = 12'h0;
    rob_1_22_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b101101))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101101))
      begin
        rob_1_22_com_1 = soc1.core.rob.rob_uop_1_22_br_mask;
        rob_1_22_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_22_com_1 = 12'h0;
        rob_1_22_uncom_1 = soc1.core.rob.rob_uop_1_22_br_mask;
      end
    end
  end

  wire [11:0] rob_1_23_com_1;
  wire [11:0] rob_1_23_uncom_1;

  always @(*)
  begin
    rob_1_23_com_1 = 12'h0;
    rob_1_23_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b101111))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b101111))
      begin
        rob_1_23_com_1 = soc1.core.rob.rob_uop_1_23_br_mask;
        rob_1_23_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_23_com_1 = 12'h0;
        rob_1_23_uncom_1 = soc1.core.rob.rob_uop_1_23_br_mask;
      end
    end
  end

  wire [11:0] rob_1_24_com_1;
  wire [11:0] rob_1_24_uncom_1;

  always @(*)
  begin
    rob_1_24_com_1 = 12'h0;
    rob_1_24_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b110001))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110001))
      begin
        rob_1_24_com_1 = soc1.core.rob.rob_uop_1_24_br_mask;
        rob_1_24_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_24_com_1 = 12'h0;
        rob_1_24_uncom_1 = soc1.core.rob.rob_uop_1_24_br_mask;
      end
    end
  end

  wire [11:0] rob_1_25_com_1;
  wire [11:0] rob_1_25_uncom_1;

  always @(*)
  begin
    rob_1_25_com_1 = 12'h0;
    rob_1_25_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b110011))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110011))
      begin
        rob_1_25_com_1 = soc1.core.rob.rob_uop_1_25_br_mask;
        rob_1_25_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_25_com_1 = 12'h0;
        rob_1_25_uncom_1 = soc1.core.rob.rob_uop_1_25_br_mask;
      end
    end
  end

  wire [11:0] rob_1_26_com_1;
  wire [11:0] rob_1_26_uncom_1;

  always @(*)
  begin
    rob_1_26_com_1 = 12'h0;
    rob_1_26_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b110101))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110101))
      begin
        rob_1_26_com_1 = soc1.core.rob.rob_uop_1_26_br_mask;
        rob_1_26_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_26_com_1 = 12'h0;
        rob_1_26_uncom_1 = soc1.core.rob.rob_uop_1_26_br_mask;
      end
    end
  end

  wire [11:0] rob_1_27_com_1;
  wire [11:0] rob_1_27_uncom_1;

  always @(*)
  begin
    rob_1_27_com_1 = 12'h0;
    rob_1_27_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b110111))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b110111))
      begin
        rob_1_27_com_1 = soc1.core.rob.rob_uop_1_27_br_mask;
        rob_1_27_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_27_com_1 = 12'h0;
        rob_1_27_uncom_1 = soc1.core.rob.rob_uop_1_27_br_mask;
      end
    end
  end

  wire [11:0] rob_1_28_com_1;
  wire [11:0] rob_1_28_uncom_1;

  always @(*)
  begin
    rob_1_28_com_1 = 12'h0;
    rob_1_28_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b111001))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111001))
      begin
        rob_1_28_com_1 = soc1.core.rob.rob_uop_1_28_br_mask;
        rob_1_28_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_28_com_1 = 12'h0;
        rob_1_28_uncom_1 = soc1.core.rob.rob_uop_1_28_br_mask;
      end
    end
  end

  wire [11:0] rob_1_29_com_1;
  wire [11:0] rob_1_29_uncom_1;

  always @(*)
  begin
    rob_1_29_com_1 = 12'h0;
    rob_1_29_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b111011))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111011))
      begin
        rob_1_29_com_1 = soc1.core.rob.rob_uop_1_29_br_mask;
        rob_1_29_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_29_com_1 = 12'h0;
        rob_1_29_uncom_1 = soc1.core.rob.rob_uop_1_29_br_mask;
      end
    end
  end

  wire [11:0] rob_1_30_com_1;
  wire [11:0] rob_1_30_uncom_1;

  always @(*)
  begin
    rob_1_30_com_1 = 12'h0;
    rob_1_30_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b111101))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111101))
      begin
        rob_1_30_com_1 = soc1.core.rob.rob_uop_1_30_br_mask;
        rob_1_30_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_30_com_1 = 12'h0;
        rob_1_30_uncom_1 = soc1.core.rob.rob_uop_1_30_br_mask;
      end
    end
  end

  wire [11:0] rob_1_31_com_1;
  wire [11:0] rob_1_31_uncom_1;

  always @(*)
  begin
    rob_1_31_com_1 = 12'h0;
    rob_1_31_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(6'b111111))
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, 6'b111111))
      begin
        rob_1_31_com_1 = soc1.core.rob.rob_uop_1_31_br_mask;
        rob_1_31_uncom_1 = 12'hfff;
      end
      else
      begin
        rob_1_31_com_1 = 12'h0;
        rob_1_31_uncom_1 = soc1.core.rob.rob_uop_1_31_br_mask;
      end
    end
  end

  wire [11:0] lsu_clr_bsy_brmask_0_com_1;
  wire [11:0] lsu_clr_bsy_brmask_0_uncom_1;

  always @(*)
  begin
    lsu_clr_bsy_brmask_0_com_1 = 12'h0;
    lsu_clr_bsy_brmask_0_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.clr_bsy_rob_idx_0) && soc1.lsu.clr_bsy_valid_0)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.clr_bsy_rob_idx_0))
      begin
        lsu_clr_bsy_brmask_0_com_1 = soc1.lsu.clr_bsy_brmask_0;
        lsu_clr_bsy_brmask_0_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_clr_bsy_brmask_0_com_1 = 12'h0;
        lsu_clr_bsy_brmask_0_uncom_1 = soc1.lsu.clr_bsy_brmask_0;
      end
    end
  end

  wire [11:0] lsu_r_xcpt_com_1;
  wire [11:0] lsu_r_xcpt_uncom_1;

  always @(*)
  begin
    lsu_r_xcpt_com_1 = 12'h0;
    lsu_r_xcpt_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(soc1.lsu.r_xcpt_uop_rob_idx) && soc1.lsu.r_xcpt_valid)
    begin
      if (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.r_xcpt_uop_rob_idx))
      begin
        lsu_r_xcpt_com_1 = soc1.lsu.r_xcpt_uop_br_mask;
        lsu_r_xcpt_uncom_1 = 12'hfff;
      end
      else
      begin
        lsu_r_xcpt_com_1 = 12'h0;
        lsu_r_xcpt_uncom_1 = soc1.lsu.r_xcpt_uop_br_mask;
      end
    end
  end

//bookkeeping buffers without explicit rob_idx
//check if loadqueue/storequeue are used and get ROB ID from ldq_idx/stq_idx

  wire [11:0] respq_uops_0_ldq_com_1;
  wire [11:0] respq_uops_0_ldq_uncom_1;

  always @(*)
  begin
    respq_uops_0_ldq_com_1 = 12'h0;
    respq_uops_0_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_0_ldq_idx]) && soc1.dcache.mshrs.respq.valids_0)
    begin
      if(soc1.dcache.mshrs.respq.uops_0_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_0_ldq_idx]))
        begin
          respq_uops_0_ldq_com_1 = soc1.dcache.mshrs.respq.uops_0_br_mask;
          respq_uops_0_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          respq_uops_0_ldq_com_1 = 12'h0;
          respq_uops_0_ldq_uncom_1 = soc1.dcache.mshrs.respq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_1_ldq_com_1;
  wire [11:0] respq_uops_1_ldq_uncom_1;

  always @(*)
  begin
    respq_uops_1_ldq_com_1 = 12'h0;
    respq_uops_1_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_1_ldq_idx]) && soc1.dcache.mshrs.respq.valids_1)
    begin
      if(soc1.dcache.mshrs.respq.uops_1_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_1_ldq_idx]))
        begin
          respq_uops_1_ldq_com_1 = soc1.dcache.mshrs.respq.uops_1_br_mask;
          respq_uops_1_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          respq_uops_1_ldq_com_1 = 12'h0;
          respq_uops_1_ldq_uncom_1 = soc1.dcache.mshrs.respq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_2_ldq_com_1;
  wire [11:0] respq_uops_2_ldq_uncom_1;

  always @(*)
  begin
    respq_uops_2_ldq_com_1 = 12'h0;
    respq_uops_2_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_2_ldq_idx]) && soc1.dcache.mshrs.respq.valids_2)
    begin
      if(soc1.dcache.mshrs.respq.uops_2_uses_ldq == 1'b1)
      begin
      if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_2_ldq_idx]))
        begin
          respq_uops_2_ldq_com_1 = soc1.dcache.mshrs.respq.uops_2_br_mask;
          respq_uops_2_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          respq_uops_2_ldq_com_1 = 12'h0;
          respq_uops_2_ldq_uncom_1 = soc1.dcache.mshrs.respq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_3_ldq_com_1;
  wire [11:0] respq_uops_3_ldq_uncom_1;

  always @(*)
  begin
    respq_uops_3_ldq_com_1 = 12'h0;
    respq_uops_3_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_3_ldq_idx]) && soc1.dcache.mshrs.respq.valids_3)
    begin
      if(soc1.dcache.mshrs.respq.uops_3_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_3_ldq_idx]))
        begin
          respq_uops_3_ldq_com_1 = soc1.dcache.mshrs.respq.uops_3_br_mask;
          respq_uops_3_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          respq_uops_3_ldq_com_1 = 12'h0;
          respq_uops_3_ldq_uncom_1 = soc1.dcache.mshrs.respq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_0_stq_com_1;
  wire [11:0] respq_uops_0_stq_uncom_1;

  always @(*)
  begin
    respq_uops_0_stq_com_1 = 12'h0;
    respq_uops_0_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_0_stq_idx]) && soc1.dcache.mshrs.respq.valids_0 && !(soc1.dcache.mshrs.respq.uops_0_uses_stq && stq_committed_1[soc1.dcache.mshrs.respq.uops_0_stq_idx]))
    begin
      if(soc1.dcache.mshrs.respq.uops_0_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_0_stq_idx]))
        begin
          respq_uops_0_stq_com_1 = soc1.dcache.mshrs.respq.uops_0_br_mask;
          respq_uops_0_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          respq_uops_0_stq_com_1 = 12'h0;
          respq_uops_0_stq_uncom_1 = soc1.dcache.mshrs.respq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_1_stq_com_1;
  wire [11:0] respq_uops_1_stq_uncom_1;

  always @(*)
  begin
    respq_uops_1_stq_com_1 = 12'h0;
    respq_uops_1_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_1_stq_idx]) && soc1.dcache.mshrs.respq.valids_1 && !(soc1.dcache.mshrs.respq.uops_1_uses_stq && stq_committed_1[soc1.dcache.mshrs.respq.uops_1_stq_idx]))
    begin
      if(soc1.dcache.mshrs.respq.uops_1_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_1_stq_idx]))
        begin
          respq_uops_1_stq_com_1 = soc1.dcache.mshrs.respq.uops_1_br_mask;
          respq_uops_1_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          respq_uops_1_stq_com_1 = 12'h0;
          respq_uops_1_stq_uncom_1 = soc1.dcache.mshrs.respq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_2_stq_com_1;
  wire [11:0] respq_uops_2_stq_uncom_1;

  always @(*)
  begin
    respq_uops_2_stq_com_1 = 12'h0;
    respq_uops_2_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_2_stq_idx]) && soc1.dcache.mshrs.respq.valids_2 && !(soc1.dcache.mshrs.respq.uops_2_uses_stq && stq_committed_1[soc1.dcache.mshrs.respq.uops_2_stq_idx]))
    begin
      if(soc1.dcache.mshrs.respq.uops_2_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_2_stq_idx]))
        begin
          respq_uops_2_stq_com_1 = soc1.dcache.mshrs.respq.uops_2_br_mask;
          respq_uops_2_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          respq_uops_2_stq_com_1 = 12'h0;
          respq_uops_2_stq_uncom_1 = soc1.dcache.mshrs.respq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_3_stq_com_1;
  wire [11:0] respq_uops_3_stq_uncom_1;

  always @(*)
  begin
    respq_uops_3_stq_com_1 = 12'h0;
    respq_uops_3_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_3_stq_idx]) && soc1.dcache.mshrs.respq.valids_3 && !(soc1.dcache.mshrs.respq.uops_3_uses_stq && stq_committed_1[soc1.dcache.mshrs.respq.uops_3_stq_idx]))
    begin
      if(soc1.dcache.mshrs.respq.uops_3_uses_stq == 1'b1)
      begin
      if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_3_stq_idx]))
        begin
          respq_uops_3_stq_com_1 = soc1.dcache.mshrs.respq.uops_3_br_mask;
          respq_uops_3_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          respq_uops_3_stq_com_1 = 12'h0;
          respq_uops_3_stq_uncom_1 = soc1.dcache.mshrs.respq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mmios_0_ldq_com_1;
  wire [11:0] mmios_0_ldq_uncom_1;

  always @(*)
  begin
    mmios_0_ldq_com_1 = 12'h0;
    mmios_0_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mmios_0.req_uop_ldq_idx]) && soc1.dcache.mshrs.mmios_0.state != 2'b0)
    begin
      if(soc1.dcache.mshrs.mmios_0.req_uop_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mmios_0.req_uop_ldq_idx]))
        begin
          mmios_0_ldq_com_1 = soc1.dcache.mshrs.mmios_0.req_uop_br_mask;
          mmios_0_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mmios_0_ldq_com_1 = 12'h0;
          mmios_0_ldq_uncom_1 = soc1.dcache.mshrs.mmios_0.req_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] mmios_0_stq_com_1;
  wire [11:0] mmios_0_stq_uncom_1;

  always @(*)
  begin
    mmios_0_stq_com_1 = 12'h0;
    mmios_0_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mmios_0.req_uop_stq_idx]) && soc1.dcache.mshrs.mmios_0.state != 2'b0)
    begin
      if((soc1.dcache.mshrs.mmios_0.req_uop_uses_stq == 1'b1) && !stq_committed_1[soc1.dcache.mshrs.mmios_0.req_uop_stq_idx])
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mmios_0.req_uop_stq_idx]))
        begin
          mmios_0_stq_com_1 = soc1.dcache.mshrs.mmios_0.req_uop_br_mask;
          mmios_0_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mmios_0_stq_com_1 = 12'h0;
          mmios_0_stq_uncom_1 = soc1.dcache.mshrs.mmios_0.req_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_0_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_0_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_0_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_0_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_0_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_0)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_0_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_0_ldq_idx]))
        begin
          mshrs_0_rpq_uops_0_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask;
          mshrs_0_rpq_uops_0_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_0_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_0_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_1_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_1_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_1_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_1_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_1_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_1)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_1_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_1_ldq_idx]))
        begin
          mshrs_0_rpq_uops_1_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask;
          mshrs_0_rpq_uops_1_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_1_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_1_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_2_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_2_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_2_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_2_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_2_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_2)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_2_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_2_ldq_idx]))
        begin
          mshrs_0_rpq_uops_2_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask;
          mshrs_0_rpq_uops_2_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_2_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_2_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_3_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_3_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_3_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_3_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_3_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_3)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_3_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_3_ldq_idx]))
        begin
          mshrs_0_rpq_uops_3_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask;
          mshrs_0_rpq_uops_3_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_3_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_3_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_4_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_4_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_4_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_4_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_4_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_4)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_4_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_4_ldq_idx]))
        begin
          mshrs_0_rpq_uops_4_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask;
          mshrs_0_rpq_uops_4_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_4_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_4_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_5_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_5_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_5_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_5_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_5_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_5)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_5_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_5_ldq_idx]))
        begin
          mshrs_0_rpq_uops_5_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask;
          mshrs_0_rpq_uops_5_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_5_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_5_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_6_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_6_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_6_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_6_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_6_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_6)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_6_uses_ldq == 1'b1)
      begin
      if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_6_ldq_idx]))
        begin
          mshrs_0_rpq_uops_6_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask;
          mshrs_0_rpq_uops_6_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_6_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_6_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_7_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_7_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_7_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_7_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_7_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_7)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_7_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_7_ldq_idx]))
        begin
          mshrs_0_rpq_uops_7_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask;
          mshrs_0_rpq_uops_7_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_7_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_7_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_8_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_8_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_8_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_8_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_8_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_8)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_8_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_8_ldq_idx]))
        begin
          mshrs_0_rpq_uops_8_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask;
          mshrs_0_rpq_uops_8_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_8_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_8_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_9_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_9_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_9_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_9_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_9_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_9)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_9_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_9_ldq_idx]))
        begin
          mshrs_0_rpq_uops_9_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask;
          mshrs_0_rpq_uops_9_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_9_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_9_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_10_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_10_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_10_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_10_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_10_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_10)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_10_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_10_ldq_idx]))
        begin
          mshrs_0_rpq_uops_10_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask;
          mshrs_0_rpq_uops_10_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_10_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_10_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_11_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_11_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_11_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_11_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_11_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_11)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_11_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_11_ldq_idx]))
        begin
          mshrs_0_rpq_uops_11_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask;
          mshrs_0_rpq_uops_11_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_11_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_11_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_12_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_12_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_12_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_12_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_12_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_12)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_12_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_12_ldq_idx]))
        begin
          mshrs_0_rpq_uops_12_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask;
          mshrs_0_rpq_uops_12_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_12_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_12_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_13_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_13_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_13_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_13_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_13_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_13)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_13_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_13_ldq_idx]))
        begin
          mshrs_0_rpq_uops_13_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask;
          mshrs_0_rpq_uops_13_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_13_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_13_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_14_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_14_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_14_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_14_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_14_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_14)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_14_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_14_ldq_idx]))
        begin
          mshrs_0_rpq_uops_14_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask;
          mshrs_0_rpq_uops_14_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_14_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_14_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_15_ldq_com_1;
  wire [11:0] mshrs_0_rpq_uops_15_ldq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_15_ldq_com_1 = 12'h0;
    mshrs_0_rpq_uops_15_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_15_ldq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_15)
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_15_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_15_ldq_idx]))
        begin
          mshrs_0_rpq_uops_15_ldq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask;
          mshrs_0_rpq_uops_15_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_15_ldq_com_1 = 12'h0;
          mshrs_0_rpq_uops_15_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask;
        end
      end
    end
  end


  wire [11:0] mshrs_0_rpq_uops_0_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_0_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_0_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_0_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_0 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_0_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx]))
        begin
          mshrs_0_rpq_uops_0_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask;
          mshrs_0_rpq_uops_0_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_0_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_0_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_1_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_1_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_1_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_1_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_1 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_1_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx]))
        begin
          mshrs_0_rpq_uops_1_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask;
          mshrs_0_rpq_uops_1_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_1_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_1_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_2_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_2_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_2_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_2_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_2 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_2_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx]))
        begin
          mshrs_0_rpq_uops_2_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask;
          mshrs_0_rpq_uops_2_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_2_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_2_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_3_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_3_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_3_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_3_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_3 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_3_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx]))
        begin
          mshrs_0_rpq_uops_3_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask;
          mshrs_0_rpq_uops_3_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_3_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_3_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_4_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_4_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_4_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_4_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_4 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_4_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx]))
        begin
          mshrs_0_rpq_uops_4_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask;
          mshrs_0_rpq_uops_4_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_4_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_4_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_5_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_5_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_5_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_5_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_5 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_5_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx]))
        begin
          mshrs_0_rpq_uops_5_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask;
          mshrs_0_rpq_uops_5_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_5_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_5_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_6_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_6_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_6_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_6_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_6 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_6_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx]))
        begin
          mshrs_0_rpq_uops_6_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask;
          mshrs_0_rpq_uops_6_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_6_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_6_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_7_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_7_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_7_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_7_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_7 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_7_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx]))
        begin
          mshrs_0_rpq_uops_7_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask;
          mshrs_0_rpq_uops_7_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_7_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_7_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_8_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_8_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_8_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_8_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_8 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_8_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx]))
        begin
          mshrs_0_rpq_uops_8_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask;
          mshrs_0_rpq_uops_8_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_8_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_8_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_9_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_9_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_9_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_9_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_9 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_9_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx]))
        begin
          mshrs_0_rpq_uops_9_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask;
          mshrs_0_rpq_uops_9_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_9_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_9_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_10_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_10_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_10_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_10_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_10 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_10_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx]))
        begin
          mshrs_0_rpq_uops_10_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask;
          mshrs_0_rpq_uops_10_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_10_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_10_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_11_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_11_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_11_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_11_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_11 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_11_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx]))
        begin
          mshrs_0_rpq_uops_11_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask;
          mshrs_0_rpq_uops_11_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_11_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_11_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_12_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_12_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_12_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_12_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_12 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_12_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx]))
        begin
          mshrs_0_rpq_uops_12_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask;
          mshrs_0_rpq_uops_12_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_12_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_12_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_13_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_13_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_13_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_13_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_13 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_13_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx]))
        begin
          mshrs_0_rpq_uops_13_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask;
          mshrs_0_rpq_uops_13_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_13_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_13_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_14_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_14_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_14_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_14_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_14 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_14_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx]))
        begin
          mshrs_0_rpq_uops_14_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask;
          mshrs_0_rpq_uops_14_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_14_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_14_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_15_stq_com_1;
  wire [11:0] mshrs_0_rpq_uops_15_stq_uncom_1;

  always @(*)
  begin
    mshrs_0_rpq_uops_15_stq_com_1 = 12'h0;
    mshrs_0_rpq_uops_15_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx]) && soc1.dcache.mshrs.mshrs_0.rpq.valids_15 && !stq_committed_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_0.rpq.uops_15_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx]))
        begin
          mshrs_0_rpq_uops_15_stq_com_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask;
          mshrs_0_rpq_uops_15_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_15_stq_com_1 = 12'h0;
          mshrs_0_rpq_uops_15_stq_uncom_1 = soc1.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_0_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_0_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_0_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_0_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_0_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_0)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_0_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_0_ldq_idx]))
        begin
          mshrs_1_rpq_uops_0_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask;
          mshrs_1_rpq_uops_0_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_0_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_0_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_1_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_1_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_1_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_1_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_1_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_1)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_1_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_1_ldq_idx]))
        begin
          mshrs_1_rpq_uops_1_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask;
          mshrs_1_rpq_uops_1_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_0_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_0_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_2_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_2_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_2_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_2_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_2_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_2)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_2_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_2_ldq_idx]))
        begin
          mshrs_1_rpq_uops_2_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask;
          mshrs_1_rpq_uops_2_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_2_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_2_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_3_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_3_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_3_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_3_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_3_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_3)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_3_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_3_ldq_idx]))
        begin
          mshrs_1_rpq_uops_3_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask;
          mshrs_1_rpq_uops_3_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_3_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_3_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_4_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_4_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_4_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_4_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_4_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_4)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_4_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_4_ldq_idx]))
        begin
          mshrs_1_rpq_uops_4_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask;
          mshrs_1_rpq_uops_4_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_4_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_4_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_5_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_5_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_5_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_5_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_5_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_5)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_5_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_5_ldq_idx]))
        begin
          mshrs_1_rpq_uops_5_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask;
          mshrs_1_rpq_uops_5_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_5_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_5_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_6_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_6_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_6_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_6_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_6_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_6)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_6_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_6_ldq_idx]))
        begin
          mshrs_1_rpq_uops_6_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask;
          mshrs_1_rpq_uops_6_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_6_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_6_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_7_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_7_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_7_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_7_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_7_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_7)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_7_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_7_ldq_idx]))
        begin
          mshrs_1_rpq_uops_7_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask;
          mshrs_1_rpq_uops_7_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_7_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_7_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_8_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_8_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_8_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_8_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_8_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_8)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_8_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_8_ldq_idx]))
        begin
          mshrs_1_rpq_uops_8_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask;
          mshrs_1_rpq_uops_8_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_8_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_8_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_9_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_9_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_9_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_9_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_9_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_9)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_9_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_9_ldq_idx]))
        begin
          mshrs_1_rpq_uops_9_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask;
          mshrs_1_rpq_uops_9_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_9_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_9_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_10_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_10_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_10_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_10_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_10_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_10)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_10_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_10_ldq_idx]))
        begin
          mshrs_1_rpq_uops_10_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask;
          mshrs_1_rpq_uops_10_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_10_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_10_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_11_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_11_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_11_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_11_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_11_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_11)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_11_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_11_ldq_idx]))
        begin
          mshrs_1_rpq_uops_11_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask;
          mshrs_1_rpq_uops_11_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_11_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_11_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_12_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_12_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_12_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_12_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_12_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_12)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_12_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_12_ldq_idx]))
        begin
          mshrs_1_rpq_uops_12_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask;
          mshrs_1_rpq_uops_12_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_12_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_12_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_13_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_13_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_13_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_13_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_13_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_13)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_13_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_13_ldq_idx]))
        begin
          mshrs_1_rpq_uops_13_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask;
          mshrs_1_rpq_uops_13_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_13_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_13_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_14_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_14_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_14_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_14_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_14_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_14)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_14_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_14_ldq_idx]))
        begin
          mshrs_1_rpq_uops_14_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask;
          mshrs_1_rpq_uops_14_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_14_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_14_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_15_ldq_com_1;
  wire [11:0] mshrs_1_rpq_uops_15_ldq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_15_ldq_com_1 = 12'h0;
    mshrs_1_rpq_uops_15_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_15_ldq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_15)
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_15_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_15_ldq_idx]))
        begin
          mshrs_1_rpq_uops_15_ldq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask;
          mshrs_1_rpq_uops_15_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_15_ldq_com_1 = 12'h0;
          mshrs_1_rpq_uops_15_ldq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask;
        end
      end
    end
  end


  wire [11:0] mshrs_1_rpq_uops_0_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_0_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_0_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_0_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_0 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_0_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx]))
        begin
          mshrs_1_rpq_uops_0_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask;
          mshrs_1_rpq_uops_0_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_0_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_0_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_1_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_1_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_1_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_1_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_1 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_1_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx]))
        begin
          mshrs_1_rpq_uops_1_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask;
          mshrs_1_rpq_uops_1_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_0_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_0_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_2_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_2_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_2_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_2_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_2 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_2_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx]))
        begin
          mshrs_1_rpq_uops_2_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask;
          mshrs_1_rpq_uops_2_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_2_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_2_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_3_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_3_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_3_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_3_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_3 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_3_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx]))
        begin
          mshrs_1_rpq_uops_3_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask;
          mshrs_1_rpq_uops_3_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_3_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_3_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_4_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_4_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_4_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_4_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_4 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_4_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx]))
        begin
          mshrs_1_rpq_uops_4_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask;
          mshrs_1_rpq_uops_4_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_4_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_4_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_5_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_5_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_5_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_5_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_5 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_5_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx]))
        begin
          mshrs_1_rpq_uops_5_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask;
          mshrs_1_rpq_uops_5_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_5_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_5_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_6_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_6_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_6_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_6_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_6 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_6_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx]))
        begin
          mshrs_1_rpq_uops_6_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask;
          mshrs_1_rpq_uops_6_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_6_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_6_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_7_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_7_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_7_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_7_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_7 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_7_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx]))
        begin
          mshrs_1_rpq_uops_7_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask;
          mshrs_1_rpq_uops_7_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_7_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_7_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_8_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_8_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_8_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_8_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_8 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_8_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx]))
        begin
          mshrs_1_rpq_uops_8_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask;
          mshrs_1_rpq_uops_8_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_8_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_8_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_9_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_9_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_9_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_9_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_9 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_9_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx]))
        begin
          mshrs_1_rpq_uops_9_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask;
          mshrs_1_rpq_uops_9_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_9_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_9_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_10_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_10_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_10_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_10_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_10 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_10_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx]))
        begin
          mshrs_1_rpq_uops_10_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask;
          mshrs_1_rpq_uops_10_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_10_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_10_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_11_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_11_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_11_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_11_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_11 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_11_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx]))
        begin
          mshrs_1_rpq_uops_11_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask;
          mshrs_1_rpq_uops_11_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_11_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_11_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_12_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_12_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_12_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_12_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_12 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_12_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx]))
        begin
          mshrs_1_rpq_uops_12_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask;
          mshrs_1_rpq_uops_12_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_12_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_12_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_13_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_13_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_13_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_13_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_13 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_13_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx]))
        begin
          mshrs_1_rpq_uops_13_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask;
          mshrs_1_rpq_uops_13_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_13_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_13_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_14_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_14_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_14_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_14_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_14 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_14_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx]))
        begin
          mshrs_1_rpq_uops_14_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask;
          mshrs_1_rpq_uops_14_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_14_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_14_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_15_stq_com_1;
  wire [11:0] mshrs_1_rpq_uops_15_stq_uncom_1;

  always @(*)
  begin
    mshrs_1_rpq_uops_15_stq_com_1 = 12'h0;
    mshrs_1_rpq_uops_15_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx]) && soc1.dcache.mshrs.mshrs_1.rpq.valids_15 && !stq_committed_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx])
    begin
      if(soc1.dcache.mshrs.mshrs_1.rpq.uops_15_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx]))
        begin
          mshrs_1_rpq_uops_15_stq_com_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask;
          mshrs_1_rpq_uops_15_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_15_stq_com_1 = 12'h0;
          mshrs_1_rpq_uops_15_stq_uncom_1 = soc1.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask;
        end
      end
    end
  end

  wire [11:0] dcache_s1_req_ldq_com_1;
  wire [11:0] dcache_s1_req_ldq_uncom_1;

  always @(*)
  begin
    dcache_s1_req_ldq_com_1 = 12'h0;
    dcache_s1_req_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.s1_req_0_uop_ldq_idx]) /*&& soc1.dcache.s1_valid_0*/)
    begin
      if(soc1.dcache.s1_req_0_uop_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.s1_req_0_uop_ldq_idx]))
        begin
          dcache_s1_req_ldq_com_1 = soc1.dcache.s1_req_0_uop_br_mask;
          dcache_s1_req_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          dcache_s1_req_ldq_com_1 = 12'h0;
          dcache_s1_req_ldq_uncom_1 = soc1.dcache.s1_req_0_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] dcache_s1_req_stq_com_1;
  wire [11:0] dcache_s1_req_stq_uncom_1;

  always @(*)
  begin
    dcache_s1_req_stq_com_1 = 12'h0;
    dcache_s1_req_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.s1_req_0_uop_stq_idx]) && /*soc1.dcache.s1_valid_0 &&*/ !stq_committed_1[soc1.dcache.s1_req_0_uop_stq_idx])
    begin
      if(soc1.dcache.s1_req_0_uop_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.s1_req_0_uop_stq_idx]))
        begin
          dcache_s1_req_stq_com_1 = soc1.dcache.s1_req_0_uop_br_mask;
          dcache_s1_req_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          dcache_s1_req_stq_com_1 = 12'h0;
          dcache_s1_req_stq_uncom_1 = soc1.dcache.s1_req_0_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] dcache_s2_req_ldq_com_1;
  wire [11:0] dcache_s2_req_ldq_uncom_1;

  always @(*)
  begin
    dcache_s2_req_ldq_com_1 = 12'h0;
    dcache_s2_req_ldq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(ldq_rob_idx_1[soc1.dcache.s2_req_0_uop_ldq_idx]) /*&& soc1.dcache.s2_valid_0*/)
    begin
      if(soc1.dcache.s2_req_0_uop_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.dcache.s2_req_0_uop_ldq_idx]))
        begin
          dcache_s2_req_ldq_com_1 = soc1.dcache.s2_req_0_uop_br_mask;
          dcache_s2_req_ldq_uncom_1 = 12'hfff;
        end
        else
        begin
          dcache_s2_req_ldq_com_1 = 12'h0;
          dcache_s2_req_ldq_uncom_1 = soc1.dcache.s2_req_0_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] dcache_s2_req_stq_com_1;
  wire [11:0] dcache_s2_req_stq_uncom_1;

  always @(*)
  begin
    dcache_s2_req_stq_com_1 = 12'h0;
    dcache_s2_req_stq_uncom_1 = 12'hfff;
    if(isInBoundsROB_1(stq_rob_idx_1[soc1.dcache.s2_req_0_uop_stq_idx]) && /*soc1.dcache.s2_valid_0 &&*/ !stq_committed_1[soc1.dcache.s2_req_0_uop_stq_idx])
    begin
      if(soc1.dcache.s2_req_0_uop_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.dcache.s2_req_0_uop_stq_idx]))
        begin
          dcache_s2_req_stq_com_1 = soc1.dcache.s2_req_0_uop_br_mask;
          dcache_s2_req_stq_uncom_1 = 12'hfff;
        end
        else
        begin
          dcache_s2_req_stq_com_1 = 12'h0;
          dcache_s2_req_stq_uncom_1 = soc1.dcache.s2_req_0_uop_br_mask;
        end
      end
    end
  end


//*******************************************//
	wire [11:0] uncommitable_masks_1;
	wire [11:0] commitable_masks_1;

//AND all uncommittable masks
assign uncommitable_masks_1 = alu_T_2_uncom_1 &
div_r_uncom_1 & exe_reg_0_uncom_1 & exe_reg_1_uncom_1 & exe_reg_2_uncom_1 & rrd_0_uncom_1 &
rrd_1_uncom_1 & rrd_2_uncom_1 & bkq_0_uncom_1 & bkq_1_uncom_1 & bkq_2_uncom_1 &
bkq_3_uncom_1 & bkq_4_uncom_1 & alu_T_2_0_uncom_1 & alu_T_2_1_uncom_1 & alu_T_2_2_uncom_1 &
ifpu_T_2_0_uncom_1 & ifpu_T_2_1_uncom_1 & imul_T_2_0_uncom_1 & imul_T_2_1_uncom_1 &
imul_T_2_2_uncom_1 & fp_issue_slot_0_uncom_1 & fp_issue_slot_1_uncom_1 & fp_issue_slot_2_uncom_1 & fp_issue_slot_3_uncom_1 &
fp_issue_slot_4_uncom_1 & fp_issue_slot_5_uncom_1 & fp_issue_slot_6_uncom_1 & fp_issue_slot_7_uncom_1 & fp_issue_slot_8_uncom_1 &
fp_issue_slot_9_uncom_1 & fp_issue_slot_10_uncom_1 & fp_issue_slot_11_uncom_1 & fp_issue_slot_12_uncom_1 & fp_issue_slot_13_uncom_1 &
fp_issue_slot_14_uncom_1 & fp_issue_slot_15_uncom_1 & fp_bkq_0_uncom_1 & fp_bkq_1_uncom_1 & fp_bkq_2_uncom_1 &
fp_bkq_3_uncom_1 & fp_bkq_4_uncom_1 & fp_bkq_5_uncom_1 & fp_bkq_6_uncom_1 & fp_bkq_1_0_uncom_1 &
fp_bkq_1_1_uncom_1 & fp_bkq_1_2_uncom_1 & fdiv_buf_uncom_1 & fdiv_divsqrt_uncom_1 & fdiv_out_uncom_1 &
fpu_T_2_0_uncom_1 & fpu_T_2_1_uncom_1 & fpu_T_2_2_uncom_1 & fpu_T_2_3_uncom_1 & f_exe_reg_uncom_1 &
f_rrd_uncom_1 & int_issue_slot_0_uncom_1 & int_issue_slot_1_uncom_1 & int_issue_slot_2_uncom_1 & int_issue_slot_3_uncom_1 &
int_issue_slot_4_uncom_1 & int_issue_slot_5_uncom_1 & int_issue_slot_6_uncom_1 & int_issue_slot_7_uncom_1 & int_issue_slot_8_uncom_1 &
int_issue_slot_9_uncom_1 & int_issue_slot_10_uncom_1 & int_issue_slot_11_uncom_1 & int_issue_slot_12_uncom_1 & int_issue_slot_13_uncom_1 &
int_issue_slot_14_uncom_1 & int_issue_slot_15_uncom_1 & int_issue_slot_16_uncom_1 & int_issue_slot_17_uncom_1 & int_issue_slot_18_uncom_1 &
int_issue_slot_19_uncom_1 & mem_issue_slot_0_uncom_1 & mem_issue_slot_1_uncom_1 & mem_issue_slot_2_uncom_1 & mem_issue_slot_3_uncom_1 &
mem_issue_slot_4_uncom_1 & mem_issue_slot_5_uncom_1 & mem_issue_slot_6_uncom_1 & mem_issue_slot_7_uncom_1 & mem_issue_slot_8_uncom_1 &
mem_issue_slot_9_uncom_1 & mem_issue_slot_10_uncom_1 & mem_issue_slot_11_uncom_1 & lsu_ldq_0_uncom_1 & lsu_ldq_1_uncom_1 &
lsu_ldq_2_uncom_1 & lsu_ldq_3_uncom_1 & lsu_ldq_4_uncom_1 & lsu_ldq_5_uncom_1 & lsu_ldq_6_uncom_1 &
lsu_ldq_7_uncom_1 & lsu_ldq_8_uncom_1 & lsu_ldq_9_uncom_1 & lsu_ldq_10_uncom_1 & lsu_ldq_11_uncom_1 &
lsu_ldq_12_uncom_1 & lsu_ldq_13_uncom_1 & lsu_ldq_14_uncom_1 & lsu_ldq_15_uncom_1 & lsu_mem_uncom_1 &
lsu_mem_stq_uncom_1 & lsu_mem_retry_uncom_1 & lsu_mem_xcpt_uncom_1 & lsu_stdf_uncom_1 & lsu_mem_stdf_uncom_1 & lsu_stq_0_uncom_1 &
lsu_stq_1_uncom_1 & lsu_stq_2_uncom_1 & lsu_stq_3_uncom_1 & lsu_stq_4_uncom_1 & lsu_stq_5_uncom_1 &
lsu_stq_6_uncom_1 & lsu_stq_7_uncom_1 & lsu_stq_8_uncom_1 & lsu_stq_9_uncom_1 & lsu_stq_10_uncom_1 &
lsu_stq_11_uncom_1 & lsu_stq_12_uncom_1 & lsu_stq_13_uncom_1 & lsu_stq_14_uncom_1 & lsu_stq_15_uncom_1 &
rob__0_uncom_1 & rob__1_uncom_1 & rob__2_uncom_1 & rob__3_uncom_1 & rob__4_uncom_1 &
rob__5_uncom_1 & rob__6_uncom_1 & rob__7_uncom_1 & rob__8_uncom_1 & rob__9_uncom_1 &
rob__10_uncom_1 & rob__11_uncom_1 & rob__12_uncom_1 & rob__13_uncom_1 & rob__14_uncom_1 &
rob__15_uncom_1 & rob__16_uncom_1 & rob__17_uncom_1 & rob__18_uncom_1 & rob__19_uncom_1 &
rob__20_uncom_1 & rob__21_uncom_1 & rob__22_uncom_1 & rob__23_uncom_1 & rob__24_uncom_1 &
rob__25_uncom_1 & rob__26_uncom_1 & rob__27_uncom_1 & rob__28_uncom_1 & rob__29_uncom_1 &
rob__30_uncom_1 & rob__31_uncom_1 & rob_1_0_uncom_1 & rob_1_1_uncom_1 & rob_1_2_uncom_1 &
rob_1_3_uncom_1 & rob_1_4_uncom_1 & rob_1_5_uncom_1 & rob_1_6_uncom_1 & rob_1_7_uncom_1 &
rob_1_8_uncom_1 & rob_1_9_uncom_1 & rob_1_10_uncom_1 & rob_1_11_uncom_1 & rob_1_12_uncom_1 &
rob_1_13_uncom_1 & rob_1_14_uncom_1 & rob_1_15_uncom_1 & rob_1_16_uncom_1 & rob_1_17_uncom_1 &
rob_1_18_uncom_1 & rob_1_19_uncom_1 & rob_1_20_uncom_1 & rob_1_21_uncom_1 & rob_1_22_uncom_1 &
rob_1_23_uncom_1 & rob_1_24_uncom_1 & rob_1_25_uncom_1 & rob_1_26_uncom_1 & rob_1_27_uncom_1 &
rob_1_28_uncom_1 & rob_1_29_uncom_1 & rob_1_30_uncom_1 & rob_1_31_uncom_1 &
lsu_clr_bsy_brmask_0_uncom_1 &
respq_uops_0_ldq_uncom_1 & respq_uops_1_ldq_uncom_1 & respq_uops_2_ldq_uncom_1 & respq_uops_3_ldq_uncom_1 &
respq_uops_0_stq_uncom_1 & respq_uops_1_stq_uncom_1 & respq_uops_2_stq_uncom_1 & respq_uops_3_stq_uncom_1 &
mmios_0_ldq_uncom_1 & mmios_0_stq_uncom_1 &
mshrs_0_rpq_uops_0_ldq_uncom_1 & mshrs_0_rpq_uops_1_ldq_uncom_1 & mshrs_0_rpq_uops_2_ldq_uncom_1 & mshrs_0_rpq_uops_3_ldq_uncom_1 &
mshrs_0_rpq_uops_4_ldq_uncom_1 & mshrs_0_rpq_uops_5_ldq_uncom_1 & mshrs_0_rpq_uops_6_ldq_uncom_1 & mshrs_0_rpq_uops_7_ldq_uncom_1 &
mshrs_0_rpq_uops_8_ldq_uncom_1 & mshrs_0_rpq_uops_9_ldq_uncom_1 & mshrs_0_rpq_uops_10_ldq_uncom_1 & mshrs_0_rpq_uops_11_ldq_uncom_1 &
mshrs_0_rpq_uops_12_ldq_uncom_1 & mshrs_0_rpq_uops_13_ldq_uncom_1 & mshrs_0_rpq_uops_14_ldq_uncom_1 & mshrs_0_rpq_uops_15_ldq_uncom_1 &/*
mshrs_0_rpq_uops_0_stq_uncom_1 & mshrs_0_rpq_uops_1_stq_uncom_1 & mshrs_0_rpq_uops_2_stq_uncom_1 & mshrs_0_rpq_uops_3_stq_uncom_1 &
mshrs_0_rpq_uops_4_stq_uncom_1 & mshrs_0_rpq_uops_5_stq_uncom_1 & mshrs_0_rpq_uops_6_stq_uncom_1 & mshrs_0_rpq_uops_7_stq_uncom_1 &
mshrs_0_rpq_uops_8_stq_uncom_1 & mshrs_0_rpq_uops_9_stq_uncom_1 & mshrs_0_rpq_uops_10_stq_uncom_1 & mshrs_0_rpq_uops_11_stq_uncom_1 &
mshrs_0_rpq_uops_12_stq_uncom_1 & mshrs_0_rpq_uops_13_stq_uncom_1 & mshrs_0_rpq_uops_14_stq_uncom_1 & mshrs_0_rpq_uops_15_stq_uncom_1 &*/
mshrs_1_rpq_uops_0_ldq_uncom_1 & mshrs_1_rpq_uops_1_ldq_uncom_1 & mshrs_1_rpq_uops_2_ldq_uncom_1 & mshrs_1_rpq_uops_3_ldq_uncom_1 &
mshrs_1_rpq_uops_4_ldq_uncom_1 & mshrs_1_rpq_uops_5_ldq_uncom_1 & mshrs_1_rpq_uops_6_ldq_uncom_1 & mshrs_1_rpq_uops_7_ldq_uncom_1 &
mshrs_1_rpq_uops_8_ldq_uncom_1 & mshrs_1_rpq_uops_9_ldq_uncom_1 & mshrs_1_rpq_uops_10_ldq_uncom_1 & mshrs_1_rpq_uops_11_ldq_uncom_1 &
mshrs_1_rpq_uops_12_ldq_uncom_1 & mshrs_1_rpq_uops_13_ldq_uncom_1 & mshrs_1_rpq_uops_14_ldq_uncom_1 & mshrs_1_rpq_uops_15_ldq_uncom_1 &/*
mshrs_1_rpq_uops_0_stq_uncom_1 & mshrs_1_rpq_uops_1_stq_uncom_1 & mshrs_1_rpq_uops_2_stq_uncom_1 & mshrs_1_rpq_uops_3_stq_uncom_1 &
mshrs_1_rpq_uops_4_stq_uncom_1 & mshrs_1_rpq_uops_5_stq_uncom_1 & mshrs_1_rpq_uops_6_stq_uncom_1 & mshrs_1_rpq_uops_7_stq_uncom_1 &
mshrs_1_rpq_uops_8_stq_uncom_1 & mshrs_1_rpq_uops_9_stq_uncom_1 & mshrs_1_rpq_uops_10_stq_uncom_1 & mshrs_1_rpq_uops_11_stq_uncom_1 &
mshrs_1_rpq_uops_12_stq_uncom_1 & mshrs_1_rpq_uops_13_stq_uncom_1 & mshrs_1_rpq_uops_14_stq_uncom_1 & mshrs_1_rpq_uops_15_stq_uncom_1 &*/
lsu_r_xcpt_uncom_1 & dcache_s1_req_ldq_uncom_1 & /*dcache_s1_req_stq_uncom_1 &*/ dcache_s2_req_ldq_uncom_1 /*& dcache_s2_req_stq_uncom_1*/;

//OR all committable masks
assign commitable_masks_1 = root_br_mask | alu_T_2_com_1 |
div_r_com_1 | exe_reg_0_com_1 | exe_reg_1_com_1 | exe_reg_2_com_1 | rrd_0_com_1 |
rrd_1_com_1 | rrd_2_com_1 | bkq_0_com_1 | bkq_1_com_1 | bkq_2_com_1 |
bkq_3_com_1 | bkq_4_com_1 | alu_T_2_0_com_1 | alu_T_2_1_com_1 | alu_T_2_2_com_1 |
ifpu_T_2_0_com_1 | ifpu_T_2_1_com_1 | imul_T_2_0_com_1 | imul_T_2_1_com_1 |
imul_T_2_2_com_1 | fp_issue_slot_0_com_1 | fp_issue_slot_1_com_1 | fp_issue_slot_2_com_1 | fp_issue_slot_3_com_1 |
fp_issue_slot_4_com_1 | fp_issue_slot_5_com_1 | fp_issue_slot_6_com_1 | fp_issue_slot_7_com_1 | fp_issue_slot_8_com_1 |
fp_issue_slot_9_com_1 | fp_issue_slot_10_com_1 | fp_issue_slot_11_com_1 | fp_issue_slot_12_com_1 | fp_issue_slot_13_com_1 |
fp_issue_slot_14_com_1 | fp_issue_slot_15_com_1 | fp_bkq_0_com_1 | fp_bkq_1_com_1 | fp_bkq_2_com_1 |
fp_bkq_3_com_1 | fp_bkq_4_com_1 | fp_bkq_5_com_1 | fp_bkq_6_com_1 | fp_bkq_1_0_com_1 |
fp_bkq_1_1_com_1 | fp_bkq_1_2_com_1 | fdiv_buf_com_1 | fdiv_divsqrt_com_1 | fdiv_out_com_1 |
fpu_T_2_0_com_1 | fpu_T_2_1_com_1 | fpu_T_2_2_com_1 | fpu_T_2_3_com_1 | f_exe_reg_com_1 |
f_rrd_com_1 | int_issue_slot_0_com_1 | int_issue_slot_1_com_1 | int_issue_slot_2_com_1 | int_issue_slot_3_com_1 |
int_issue_slot_4_com_1 | int_issue_slot_5_com_1 | int_issue_slot_6_com_1 | int_issue_slot_7_com_1 | int_issue_slot_8_com_1 |
int_issue_slot_9_com_1 | int_issue_slot_10_com_1 | int_issue_slot_11_com_1 | int_issue_slot_12_com_1 | int_issue_slot_13_com_1 |
int_issue_slot_14_com_1 | int_issue_slot_15_com_1 | int_issue_slot_16_com_1 | int_issue_slot_17_com_1 | int_issue_slot_18_com_1 |
int_issue_slot_19_com_1 | mem_issue_slot_0_com_1 | mem_issue_slot_1_com_1 | mem_issue_slot_2_com_1 | mem_issue_slot_3_com_1 |
mem_issue_slot_4_com_1 | mem_issue_slot_5_com_1 | mem_issue_slot_6_com_1 | mem_issue_slot_7_com_1 | mem_issue_slot_8_com_1 |
mem_issue_slot_9_com_1 | mem_issue_slot_10_com_1 | mem_issue_slot_11_com_1 | lsu_ldq_0_com_1 | lsu_ldq_1_com_1 |
lsu_ldq_2_com_1 | lsu_ldq_3_com_1 | lsu_ldq_4_com_1 | lsu_ldq_5_com_1 | lsu_ldq_6_com_1 |
lsu_ldq_7_com_1 | lsu_ldq_8_com_1 | lsu_ldq_9_com_1 | lsu_ldq_10_com_1 | lsu_ldq_11_com_1 |
lsu_ldq_12_com_1 | lsu_ldq_13_com_1 | lsu_ldq_14_com_1 | lsu_ldq_15_com_1 | lsu_mem_com_1 |
lsu_mem_stq_com_1 | lsu_mem_retry_com_1 | lsu_mem_xcpt_com_1 | lsu_stdf_com_1 | lsu_mem_stdf_com_1 | lsu_stq_0_com_1 |
lsu_stq_1_com_1 | lsu_stq_2_com_1 | lsu_stq_3_com_1 | lsu_stq_4_com_1 | lsu_stq_5_com_1 |
lsu_stq_6_com_1 | lsu_stq_7_com_1 | lsu_stq_8_com_1 | lsu_stq_9_com_1 | lsu_stq_10_com_1 |
lsu_stq_11_com_1 | lsu_stq_12_com_1 | lsu_stq_13_com_1 | lsu_stq_14_com_1 | lsu_stq_15_com_1 |
rob__0_com_1 | rob__1_com_1 | rob__2_com_1 | rob__3_com_1 | rob__4_com_1 |
rob__5_com_1 | rob__6_com_1 | rob__7_com_1 | rob__8_com_1 | rob__9_com_1 |
rob__10_com_1 | rob__11_com_1 | rob__12_com_1 | rob__13_com_1 | rob__14_com_1 |
rob__15_com_1 | rob__16_com_1 | rob__17_com_1 | rob__18_com_1 | rob__19_com_1 |
rob__20_com_1 | rob__21_com_1 | rob__22_com_1 | rob__23_com_1 | rob__24_com_1 |
rob__25_com_1 | rob__26_com_1 | rob__27_com_1 | rob__28_com_1 | rob__29_com_1 |
rob__30_com_1 | rob__31_com_1 | rob_1_0_com_1 | rob_1_1_com_1 | rob_1_2_com_1 |
rob_1_3_com_1 | rob_1_4_com_1 | rob_1_5_com_1 | rob_1_6_com_1 | rob_1_7_com_1 |
rob_1_8_com_1 | rob_1_9_com_1 | rob_1_10_com_1 | rob_1_11_com_1 | rob_1_12_com_1 |
rob_1_13_com_1 | rob_1_14_com_1 | rob_1_15_com_1 | rob_1_16_com_1 | rob_1_17_com_1 |
rob_1_18_com_1 | rob_1_19_com_1 | rob_1_20_com_1 | rob_1_21_com_1 | rob_1_22_com_1 |
rob_1_23_com_1 | rob_1_24_com_1 | rob_1_25_com_1 | rob_1_26_com_1 | rob_1_27_com_1 |
rob_1_28_com_1 | rob_1_29_com_1 | rob_1_30_com_1 | rob_1_31_com_1 |
lsu_clr_bsy_brmask_0_com_1 |
respq_uops_0_ldq_com_1 | respq_uops_1_ldq_com_1 | respq_uops_2_ldq_com_1 | respq_uops_3_ldq_com_1 |
respq_uops_0_stq_com_1 | respq_uops_1_stq_com_1 | respq_uops_2_stq_com_1 | respq_uops_3_stq_com_1 |
mmios_0_ldq_com_1 | mmios_0_stq_com_1 |
mshrs_0_rpq_uops_0_ldq_com_1 | mshrs_0_rpq_uops_1_ldq_com_1 | mshrs_0_rpq_uops_2_ldq_com_1 | mshrs_0_rpq_uops_3_ldq_com_1 |
mshrs_0_rpq_uops_4_ldq_com_1 | mshrs_0_rpq_uops_5_ldq_com_1 | mshrs_0_rpq_uops_6_ldq_com_1 | mshrs_0_rpq_uops_7_ldq_com_1 |
mshrs_0_rpq_uops_8_ldq_com_1 | mshrs_0_rpq_uops_9_ldq_com_1 | mshrs_0_rpq_uops_10_ldq_com_1 | mshrs_0_rpq_uops_11_ldq_com_1 |
mshrs_0_rpq_uops_12_ldq_com_1 | mshrs_0_rpq_uops_13_ldq_com_1 | mshrs_0_rpq_uops_14_ldq_com_1 | mshrs_0_rpq_uops_15_ldq_com_1 |/*
mshrs_0_rpq_uops_0_stq_com_1 | mshrs_0_rpq_uops_1_stq_com_1 | mshrs_0_rpq_uops_2_stq_com_1 | mshrs_0_rpq_uops_3_stq_com_1 |
mshrs_0_rpq_uops_4_stq_com_1 | mshrs_0_rpq_uops_5_stq_com_1 | mshrs_0_rpq_uops_6_stq_com_1 | mshrs_0_rpq_uops_7_stq_com_1 |
mshrs_0_rpq_uops_8_stq_com_1 | mshrs_0_rpq_uops_9_stq_com_1 | mshrs_0_rpq_uops_10_stq_com_1 | mshrs_0_rpq_uops_11_stq_com_1 |
mshrs_0_rpq_uops_12_stq_com_1 | mshrs_0_rpq_uops_13_stq_com_1 | mshrs_0_rpq_uops_14_stq_com_1 | mshrs_0_rpq_uops_15_stq_com_1 |*/
mshrs_1_rpq_uops_0_ldq_com_1 | mshrs_1_rpq_uops_1_ldq_com_1 | mshrs_1_rpq_uops_2_ldq_com_1 | mshrs_1_rpq_uops_3_ldq_com_1 |
mshrs_1_rpq_uops_4_ldq_com_1 | mshrs_1_rpq_uops_5_ldq_com_1 | mshrs_1_rpq_uops_6_ldq_com_1 | mshrs_1_rpq_uops_7_ldq_com_1 |
mshrs_1_rpq_uops_8_ldq_com_1 | mshrs_1_rpq_uops_9_ldq_com_1 | mshrs_1_rpq_uops_10_ldq_com_1 | mshrs_1_rpq_uops_11_ldq_com_1 |
mshrs_1_rpq_uops_12_ldq_com_1 | mshrs_1_rpq_uops_13_ldq_com_1 | mshrs_1_rpq_uops_14_ldq_com_1 | mshrs_1_rpq_uops_15_ldq_com_1 |/*
mshrs_1_rpq_uops_0_stq_com_1 | mshrs_1_rpq_uops_1_stq_com_1 | mshrs_1_rpq_uops_2_stq_com_1 | mshrs_1_rpq_uops_3_stq_com_1 |
mshrs_1_rpq_uops_4_stq_com_1 | mshrs_1_rpq_uops_5_stq_com_1 | mshrs_1_rpq_uops_6_stq_com_1 | mshrs_1_rpq_uops_7_stq_com_1 |
mshrs_1_rpq_uops_8_stq_com_1 | mshrs_1_rpq_uops_9_stq_com_1 | mshrs_1_rpq_uops_10_stq_com_1 | mshrs_1_rpq_uops_11_stq_com_1 |
mshrs_1_rpq_uops_12_stq_com_1 | mshrs_1_rpq_uops_13_stq_com_1 | mshrs_1_rpq_uops_14_stq_com_1 | mshrs_1_rpq_uops_15_stq_com_1 |*/
lsu_r_xcpt_com_1 | dcache_s1_req_ldq_com_1 | /*dcache_s1_req_stq_com_1 |*/ dcache_s2_req_ldq_com_1 /*| dcache_s2_req_stq_com_1*/;


//***************************************//
//write one combinational process for both ME-5 and ME-6
//for every ROB slot or bookkeeping buffer:
//check if stored ROB ID is committable
//store branch mask in corresponding variable
//set the other variable to default value (12'hfff for uncommitable tags, 12'h0 for committable tags)

//Soc2
//

  wire [11:0] alu_T_2_com_2;
  wire [11:0] alu_T_2_uncom_2;

  always @(*)
  begin
    alu_T_2_com_2 = 12'h0;
    alu_T_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.csr_exe_unit.alu.r_uops_0_rob_idx) && soc2.core.csr_exe_unit.alu.r_valids_0)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.csr_exe_unit.alu.r_uops_0_rob_idx))
      begin
        alu_T_2_com_2 = soc2.core.csr_exe_unit.alu.r_uops_0_br_mask;
        alu_T_2_uncom_2 = 12'hfff;
      end
      else
      begin
        alu_T_2_com_2 = 12'h0;
        alu_T_2_uncom_2 = soc2.core.csr_exe_unit.alu.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] div_r_com_2;
  wire [11:0] div_r_uncom_2;

  always @(*)
  begin
    div_r_com_2 = 12'h0;
    div_r_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.csr_exe_unit.div.r_uop_rob_idx) && (soc2.core.csr_exe_unit.div.div.state == 3'h3))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.csr_exe_unit.div.r_uop_rob_idx))
      begin
        div_r_com_2 = soc2.core.csr_exe_unit.div.r_uop_br_mask;
        div_r_uncom_2 = 12'hfff;
      end
      else
      begin
        div_r_com_2 = 12'h0;
        div_r_uncom_2 = soc2.core.csr_exe_unit.div.r_uop_br_mask;
      end
    end
  end

  wire [11:0] exe_reg_0_com_2;
  wire [11:0] exe_reg_0_uncom_2;

  always @(*)
  begin
    exe_reg_0_com_2 = 12'h0;
    exe_reg_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.iregister_read.exe_reg_uops_0_rob_idx) && soc2.core.iregister_read.exe_reg_valids_0 && !(soc2.core.iregister_read.exe_reg_uops_0_uses_stq && stq_committed_2[soc2.core.iregister_read.exe_reg_uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.exe_reg_uops_0_rob_idx))
      begin
        exe_reg_0_com_2 = soc2.core.iregister_read.exe_reg_uops_0_br_mask;
        exe_reg_0_uncom_2 = 12'hfff;
      end
      else
      begin
        exe_reg_0_com_2 = 12'h0;
        exe_reg_0_uncom_2 = soc2.core.iregister_read.exe_reg_uops_0_br_mask;
      end
    end
  end

  wire [11:0] exe_reg_1_com_2;
  wire [11:0] exe_reg_1_uncom_2;

  always @(*)
  begin
    exe_reg_1_com_2 = 12'h0;
    exe_reg_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.iregister_read.exe_reg_uops_1_rob_idx) && soc2.core.iregister_read.exe_reg_valids_1 && !(soc2.core.iregister_read.exe_reg_uops_1_uses_stq && stq_committed_2[soc2.core.iregister_read.exe_reg_uops_1_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.exe_reg_uops_1_rob_idx))
      begin
        exe_reg_1_com_2 = soc2.core.iregister_read.exe_reg_uops_1_br_mask;
        exe_reg_1_uncom_2 = 12'hfff;
      end
      else
      begin
        exe_reg_1_com_2 = 12'h0;
        exe_reg_1_uncom_2 = soc2.core.iregister_read.exe_reg_uops_1_br_mask;
      end
    end
  end

  wire [11:0] exe_reg_2_com_2;
  wire [11:0] exe_reg_2_uncom_2;

  always @(*)
  begin
    exe_reg_2_com_2 = 12'h0;
    exe_reg_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.iregister_read.exe_reg_uops_2_rob_idx) && soc2.core.iregister_read.exe_reg_valids_2 && !(soc2.core.iregister_read.exe_reg_uops_2_uses_stq && stq_committed_2[soc2.core.iregister_read.exe_reg_uops_2_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.exe_reg_uops_2_rob_idx))
      begin
        exe_reg_2_com_2 = soc2.core.iregister_read.exe_reg_uops_2_br_mask;
        exe_reg_2_uncom_2 = 12'hfff;
      end
      else
      begin
        exe_reg_2_com_2 = 12'h0;
        exe_reg_2_uncom_2 = soc2.core.iregister_read.exe_reg_uops_2_br_mask;
      end
    end
  end

  wire [11:0] rrd_0_com_2;
  wire [11:0] rrd_0_uncom_2;

  always @(*)
  begin
    rrd_0_com_2 = 12'h0;
    rrd_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.iregister_read.rrd_uops_0_REG_rob_idx) && soc2.core.iregister_read.rrd_valids_0_REG && !(soc2.core.iregister_read.rrd_uops_0_REG_uses_stq && stq_committed_2[soc2.core.iregister_read.rrd_uops_0_REG_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.rrd_uops_0_REG_rob_idx))
      begin
        rrd_0_com_2 = soc2.core.iregister_read.rrd_uops_0_REG_br_mask;
        rrd_0_uncom_2 = 12'hfff;
      end
      else
      begin
        rrd_0_com_2 = 12'h0;
        rrd_0_uncom_2 = soc2.core.iregister_read.rrd_uops_0_REG_br_mask;
      end
    end
  end

  wire [11:0] rrd_1_com_2;
  wire [11:0] rrd_1_uncom_2;

  always @(*)
  begin
    rrd_1_com_2 = 12'h0;
    rrd_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.iregister_read.rrd_uops_1_REG_rob_idx) && soc2.core.iregister_read.rrd_valids_1_REG && !(soc2.core.iregister_read.rrd_uops_1_REG_uses_stq && stq_committed_2[soc2.core.iregister_read.rrd_uops_1_REG_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.rrd_uops_1_REG_rob_idx))
      begin
        rrd_1_com_2 = soc2.core.iregister_read.rrd_uops_1_REG_br_mask;
        rrd_1_uncom_2 = 12'hfff;
      end
      else
      begin
        rrd_1_com_2 = 12'h0;
        rrd_1_uncom_2 = soc2.core.iregister_read.rrd_uops_1_REG_br_mask;
      end
    end
  end

  wire [11:0] rrd_2_com_2;
  wire [11:0] rrd_2_uncom_2;

  always @(*)
  begin
    rrd_2_com_2 = 12'h0;
    rrd_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.iregister_read.rrd_uops_2_REG_rob_idx) && soc2.core.iregister_read.rrd_valids_2_REG && !(soc2.core.iregister_read.rrd_uops_2_REG_uses_stq && stq_committed_2[soc2.core.iregister_read.rrd_uops_2_REG_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.rrd_uops_2_REG_rob_idx))
      begin
        rrd_2_com_2 = soc2.core.iregister_read.rrd_uops_2_REG_br_mask;
        rrd_2_uncom_2 = 12'hfff;
      end
      else
      begin
        rrd_2_com_2 = 12'h0;
        rrd_2_uncom_2 = soc2.core.iregister_read.rrd_uops_2_REG_br_mask;
      end
    end
  end

  wire [11:0] bkq_0_com_2;
  wire [11:0] bkq_0_uncom_2;

  always @(*)
  begin
    bkq_0_com_2 = 12'h0;
    bkq_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.queue.uops_0_rob_idx) && soc2.core.jmp_unit.queue.valids_0 /*&& !(soc2.core.jmp_unit.queue.uops_0_uses_stq && stq_committed_2[soc2.core.jmp_unit.queue.uops_0_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.queue.uops_0_rob_idx))
      begin
        bkq_0_com_2 = soc2.core.jmp_unit.queue.uops_0_br_mask;
        bkq_0_uncom_2 = 12'hfff;
      end
      else
      begin
        bkq_0_com_2 = 12'h0;
        bkq_0_uncom_2 = soc2.core.jmp_unit.queue.uops_0_br_mask;
      end
    end
  end

  wire [11:0] bkq_1_com_2;
  wire [11:0] bkq_1_uncom_2;

  always @(*)
  begin
    bkq_1_com_2 = 12'h0;
    bkq_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.queue.uops_1_rob_idx) && soc2.core.jmp_unit.queue.valids_1 /*&& !(soc2.core.jmp_unit.queue.uops_1_uses_stq && stq_committed_2[soc2.core.jmp_unit.queue.uops_1_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.queue.uops_1_rob_idx))
      begin
        bkq_1_com_2 = soc2.core.jmp_unit.queue.uops_1_br_mask;
        bkq_1_uncom_2 = 12'hfff;
      end
      else
      begin
        bkq_1_com_2 = 12'h0;
        bkq_1_uncom_2 = soc2.core.jmp_unit.queue.uops_1_br_mask;
      end
    end
  end

  wire [11:0] bkq_2_com_2;
  wire [11:0] bkq_2_uncom_2;

  always @(*)
  begin
    bkq_2_com_2 = 12'h0;
    bkq_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.queue.uops_2_rob_idx) && soc2.core.jmp_unit.queue.valids_2 /*&& !(soc2.core.jmp_unit.queue.uops_2_uses_stq && stq_committed_2[soc2.core.jmp_unit.queue.uops_2_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.queue.uops_2_rob_idx))
      begin
        bkq_2_com_2 = soc2.core.jmp_unit.queue.uops_2_br_mask;
        bkq_2_uncom_2 = 12'hfff;
      end
      else
      begin
        bkq_2_com_2 = 12'h0;
        bkq_2_uncom_2 = soc2.core.jmp_unit.queue.uops_2_br_mask;
      end
    end
  end

  wire [11:0] bkq_3_com_2;
  wire [11:0] bkq_3_uncom_2;

  always @(*)
  begin
    bkq_3_com_2 = 12'h0;
    bkq_3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.queue.uops_3_rob_idx) && soc2.core.jmp_unit.queue.valids_3 /*&& !(soc2.core.jmp_unit.queue.uops_3_uses_stq && stq_committed_2[soc2.core.jmp_unit.queue.uops_3_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.queue.uops_3_rob_idx))
      begin
        bkq_3_com_2 = soc2.core.jmp_unit.queue.uops_3_br_mask;
        bkq_3_uncom_2 = 12'hfff;
      end
      else
      begin
        bkq_3_com_2 = 12'h0;
        bkq_3_uncom_2 = soc2.core.jmp_unit.queue.uops_3_br_mask;
      end
    end
  end

  wire [11:0] bkq_4_com_2;
  wire [11:0] bkq_4_uncom_2;

  always @(*)
  begin
    bkq_4_com_2 = 12'h0;
    bkq_4_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.queue.uops_4_rob_idx) && soc2.core.jmp_unit.queue.valids_4 /*&& !(soc2.core.jmp_unit.queue.uops_4_uses_stq && stq_committed_2[soc2.core.jmp_unit.queue.uops_4_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.queue.uops_4_rob_idx))
      begin
        bkq_4_com_2 = soc2.core.jmp_unit.queue.uops_4_br_mask;
        bkq_4_uncom_2 = 12'hfff;
      end
      else
      begin
        bkq_4_com_2 = 12'h0;
        bkq_4_uncom_2 = soc2.core.jmp_unit.queue.uops_4_br_mask;
      end
    end
  end

  wire [11:0] alu_T_2_0_com_2;
  wire [11:0] alu_T_2_0_uncom_2;

  always @(*)
  begin
    alu_T_2_0_com_2 = 12'h0;
    alu_T_2_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.alu.r_uops_0_rob_idx) && soc2.core.jmp_unit.alu.r_valids_0)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.alu.r_uops_0_rob_idx))
      begin
        alu_T_2_0_com_2 = soc2.core.jmp_unit.alu.r_uops_0_br_mask;
        alu_T_2_0_uncom_2 = 12'hfff;
      end
      else
      begin
        alu_T_2_0_com_2 = 12'h0;
        alu_T_2_0_uncom_2 = soc2.core.jmp_unit.alu.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] alu_T_2_1_com_2;
  wire [11:0] alu_T_2_1_uncom_2;

  always @(*)
  begin
    alu_T_2_1_com_2 = 12'h0;
    alu_T_2_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.alu.r_uops_1_rob_idx) && soc2.core.jmp_unit.alu.r_valids_1)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.alu.r_uops_1_rob_idx))
      begin
        alu_T_2_1_com_2 = soc2.core.jmp_unit.alu.r_uops_1_br_mask;
        alu_T_2_1_uncom_2 = 12'hfff;
      end
      else
      begin
        alu_T_2_1_com_2 = 12'h0;
        alu_T_2_1_uncom_2 = soc2.core.jmp_unit.alu.r_uops_1_br_mask;
      end
    end
  end

  wire [11:0] alu_T_2_2_com_2;
  wire [11:0] alu_T_2_2_uncom_2;

  always @(*)
  begin
    alu_T_2_2_com_2 = 12'h0;
    alu_T_2_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.alu.r_uops_2_rob_idx) && soc2.core.jmp_unit.alu.r_valids_2)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.alu.r_uops_2_rob_idx))
      begin
        alu_T_2_2_com_2 = soc2.core.jmp_unit.alu.r_uops_2_br_mask;
        alu_T_2_2_uncom_2 = 12'hfff;
      end
      else
      begin
        alu_T_2_2_com_2 = 12'h0;
        alu_T_2_2_uncom_2 = soc2.core.jmp_unit.alu.r_uops_2_br_mask;
      end
    end
  end

  wire [11:0] ifpu_T_2_0_com_2;
  wire [11:0] ifpu_T_2_0_uncom_2;

  always @(*)
  begin
    ifpu_T_2_0_com_2 = 12'h0;
    ifpu_T_2_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.ifpu.r_uops_0_rob_idx) && soc2.core.jmp_unit.ifpu.r_valids_0 /*&& !(soc2.core.jmp_unit.ifpu.r_uops_0_uses_stq && stq_committed_2[soc2.core.jmp_unit.ifpu.r_uops_0_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.ifpu.r_uops_0_rob_idx))
      begin
        ifpu_T_2_0_com_2 = soc2.core.jmp_unit.ifpu.r_uops_0_br_mask;
        ifpu_T_2_0_uncom_2 = 12'hfff;
      end
      else
      begin
        ifpu_T_2_0_com_2 = 12'h0;
        ifpu_T_2_0_uncom_2 = soc2.core.jmp_unit.ifpu.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] ifpu_T_2_1_com_2;
  wire [11:0] ifpu_T_2_1_uncom_2;

  always @(*)
  begin
    ifpu_T_2_1_com_2 = 12'h0;
    ifpu_T_2_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.ifpu.r_uops_1_rob_idx) && soc2.core.jmp_unit.ifpu.r_valids_1 /*&& !(soc2.core.jmp_unit.ifpu.r_uops_1_uses_stq && stq_committed_2[soc2.core.jmp_unit.ifpu.r_uops_1_stq_idx])*/)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.ifpu.r_uops_1_rob_idx))
      begin
        ifpu_T_2_1_com_2 = soc2.core.jmp_unit.ifpu.r_uops_1_br_mask;
        ifpu_T_2_1_uncom_2 = 12'hfff;
      end
      else
      begin
        ifpu_T_2_1_com_2 = 12'h0;
        ifpu_T_2_1_uncom_2 = soc2.core.jmp_unit.ifpu.r_uops_1_br_mask;
      end
    end
  end



  wire [11:0] imul_T_2_0_com_2;
  wire [11:0] imul_T_2_0_uncom_2;

  always @(*)
  begin
    imul_T_2_0_com_2 = 12'h0;
    imul_T_2_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.imul.r_uops_0_rob_idx) && soc2.core.jmp_unit.imul.r_valids_0)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.imul.r_uops_0_rob_idx))
      begin
        imul_T_2_0_com_2 = soc2.core.jmp_unit.imul.r_uops_0_br_mask;
        imul_T_2_0_uncom_2 = 12'hfff;
      end
      else
      begin
        imul_T_2_0_com_2 = 12'h0;
        imul_T_2_0_uncom_2 = soc2.core.jmp_unit.imul.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] imul_T_2_1_com_2;
  wire [11:0] imul_T_2_1_uncom_2;

  always @(*)
  begin
    imul_T_2_1_com_2 = 12'h0;
    imul_T_2_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.imul.r_uops_1_rob_idx) && soc2.core.jmp_unit.imul.r_valids_1)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.imul.r_uops_1_rob_idx))
      begin
        imul_T_2_1_com_2 = soc2.core.jmp_unit.imul.r_uops_1_br_mask;
        imul_T_2_1_uncom_2 = 12'hfff;
      end
      else
      begin
        imul_T_2_1_com_2 = 12'h0;
        imul_T_2_1_uncom_2 = soc2.core.jmp_unit.imul.r_uops_1_br_mask;
      end
    end
  end

  wire [11:0] imul_T_2_2_com_2;
  wire [11:0] imul_T_2_2_uncom_2;

  always @(*)
  begin
    imul_T_2_2_com_2 = 12'h0;
    imul_T_2_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.jmp_unit.imul.r_uops_2_rob_idx) && soc2.core.jmp_unit.imul.r_valids_2)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.imul.r_uops_2_rob_idx))
      begin
        imul_T_2_2_com_2 = soc2.core.jmp_unit.imul.r_uops_2_br_mask;
        imul_T_2_2_uncom_2 = 12'hfff;
      end
      else
      begin
        imul_T_2_2_com_2 = 12'h0;
        imul_T_2_2_uncom_2 = soc2.core.jmp_unit.imul.r_uops_2_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_0_com_2;
  wire [11:0] fp_issue_slot_0_uncom_2;

  always @(*)
  begin
    fp_issue_slot_0_com_2 = 12'h0;
    fp_issue_slot_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_0.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx))
      begin
        fp_issue_slot_0_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_br_mask;
        fp_issue_slot_0_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_0_com_2 = 12'h0;
        fp_issue_slot_0_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_1_com_2;
  wire [11:0] fp_issue_slot_1_uncom_2;

  always @(*)
  begin
    fp_issue_slot_1_com_2 = 12'h0;
    fp_issue_slot_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_1.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx))
      begin
        fp_issue_slot_1_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_br_mask;
        fp_issue_slot_1_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_1_com_2 = 12'h0;
        fp_issue_slot_1_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_2_com_2;
  wire [11:0] fp_issue_slot_2_uncom_2;

  always @(*)
  begin
    fp_issue_slot_2_com_2 = 12'h0;
    fp_issue_slot_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_2.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx))
      begin
        fp_issue_slot_2_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_br_mask;
        fp_issue_slot_2_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_2_com_2 = 12'h0;
        fp_issue_slot_2_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_3_com_2;
  wire [11:0] fp_issue_slot_3_uncom_2;

  always @(*)
  begin
    fp_issue_slot_3_com_2 = 12'h0;
    fp_issue_slot_3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_3.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx))
      begin
        fp_issue_slot_3_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_br_mask;
        fp_issue_slot_3_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_3_com_2 = 12'h0;
        fp_issue_slot_3_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_4_com_2;
  wire [11:0] fp_issue_slot_4_uncom_2;

  always @(*)
  begin
    fp_issue_slot_4_com_2 = 12'h0;
    fp_issue_slot_4_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_4.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx))
      begin
        fp_issue_slot_4_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_br_mask;
        fp_issue_slot_4_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_4_com_2 = 12'h0;
        fp_issue_slot_4_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_5_com_2;
  wire [11:0] fp_issue_slot_5_uncom_2;

  always @(*)
  begin
    fp_issue_slot_5_com_2 = 12'h0;
    fp_issue_slot_5_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_5.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx))
      begin
        fp_issue_slot_5_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_br_mask;
        fp_issue_slot_5_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_5_com_2 = 12'h0;
        fp_issue_slot_5_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_6_com_2;
  wire [11:0] fp_issue_slot_6_uncom_2;

  always @(*)
  begin
    fp_issue_slot_6_com_2 = 12'h0;
    fp_issue_slot_6_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_6.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx))
      begin
        fp_issue_slot_6_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_br_mask;
        fp_issue_slot_6_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_6_com_2 = 12'h0;
        fp_issue_slot_6_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_7_com_2;
  wire [11:0] fp_issue_slot_7_uncom_2;

  always @(*)
  begin
    fp_issue_slot_7_com_2 = 12'h0;
    fp_issue_slot_7_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_7.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx))
      begin
        fp_issue_slot_7_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_br_mask;
        fp_issue_slot_7_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_7_com_2 = 12'h0;
        fp_issue_slot_7_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_8_com_2;
  wire [11:0] fp_issue_slot_8_uncom_2;

  always @(*)
  begin
    fp_issue_slot_8_com_2 = 12'h0;
    fp_issue_slot_8_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_8.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx))
      begin
        fp_issue_slot_8_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_br_mask;
        fp_issue_slot_8_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_8_com_2 = 12'h0;
        fp_issue_slot_8_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_9_com_2;
  wire [11:0] fp_issue_slot_9_uncom_2;

  always @(*)
  begin
    fp_issue_slot_9_com_2 = 12'h0;
    fp_issue_slot_9_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_9.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx))
      begin
        fp_issue_slot_9_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_br_mask;
        fp_issue_slot_9_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_9_com_2 = 12'h0;
        fp_issue_slot_9_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_10_com_2;
  wire [11:0] fp_issue_slot_10_uncom_2;

  always @(*)
  begin
    fp_issue_slot_10_com_2 = 12'h0;
    fp_issue_slot_10_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_10.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx))
      begin
        fp_issue_slot_10_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_br_mask;
        fp_issue_slot_10_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_10_com_2 = 12'h0;
        fp_issue_slot_10_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_11_com_2;
  wire [11:0] fp_issue_slot_11_uncom_2;

  always @(*)
  begin
    fp_issue_slot_11_com_2 = 12'h0;
    fp_issue_slot_11_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_11.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx))
      begin
        fp_issue_slot_11_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_br_mask;
        fp_issue_slot_11_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_11_com_2 = 12'h0;
        fp_issue_slot_11_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_12_com_2;
  wire [11:0] fp_issue_slot_12_uncom_2;

  always @(*)
  begin
    fp_issue_slot_12_com_2 = 12'h0;
    fp_issue_slot_12_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_12.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx))
      begin
        fp_issue_slot_12_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_br_mask;
        fp_issue_slot_12_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_12_com_2 = 12'h0;
        fp_issue_slot_12_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_13_com_2;
  wire [11:0] fp_issue_slot_13_uncom_2;

  always @(*)
  begin
    fp_issue_slot_13_com_2 = 12'h0;
    fp_issue_slot_13_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_13.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx))
      begin
        fp_issue_slot_13_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_br_mask;
        fp_issue_slot_13_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_13_com_2 = 12'h0;
        fp_issue_slot_13_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_14_com_2;
  wire [11:0] fp_issue_slot_14_uncom_2;

  always @(*)
  begin
    fp_issue_slot_14_com_2 = 12'h0;
    fp_issue_slot_14_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_14.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx))
      begin
        fp_issue_slot_14_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_br_mask;
        fp_issue_slot_14_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_14_com_2 = 12'h0;
        fp_issue_slot_14_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_issue_slot_15_com_2;
  wire [11:0] fp_issue_slot_15_uncom_2;

  always @(*)
  begin
    fp_issue_slot_15_com_2 = 12'h0;
    fp_issue_slot_15_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx) && soc2.core.fp_pipeline.fp_issue_unit.slots_15.io_valid && !(soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx))
      begin
        fp_issue_slot_15_com_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_br_mask;
        fp_issue_slot_15_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_issue_slot_15_com_2 = 12'h0;
        fp_issue_slot_15_uncom_2 = soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_0_com_2;
  wire [11:0] fp_bkq_0_uncom_2;

  always @(*)
  begin
    fp_bkq_0_com_2 = 12'h0;
    fp_bkq_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.queue.valids_0 && !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx))
      begin
        fp_bkq_0_com_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_br_mask;
        fp_bkq_0_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_0_com_2 = 12'h0;
        fp_bkq_0_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_1_com_2;
  wire [11:0] fp_bkq_1_uncom_2;

  always @(*)
  begin
    fp_bkq_1_com_2 = 12'h0;
    fp_bkq_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.queue.valids_1 && !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx))
      begin
        fp_bkq_1_com_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_br_mask;
        fp_bkq_1_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_1_com_2 = 12'h0;
        fp_bkq_1_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_2_com_2;
  wire [11:0] fp_bkq_2_uncom_2;

  always @(*)
  begin
    fp_bkq_2_com_2 = 12'h0;
    fp_bkq_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.queue.valids_2 && !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx))
      begin
        fp_bkq_2_com_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_br_mask;
        fp_bkq_2_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_2_com_2 = 12'h0;
        fp_bkq_2_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_3_com_2;
  wire [11:0] fp_bkq_3_uncom_2;

  always @(*)
  begin
    fp_bkq_3_com_2 = 12'h0;
    fp_bkq_3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.queue.valids_3 && !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx))
      begin
        fp_bkq_3_com_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_br_mask;
        fp_bkq_3_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_3_com_2 = 12'h0;
        fp_bkq_3_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_4_com_2;
  wire [11:0] fp_bkq_4_uncom_2;

  always @(*)
  begin
    fp_bkq_4_com_2 = 12'h0;
    fp_bkq_4_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.queue.valids_4 && !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx))
      begin
        fp_bkq_4_com_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_br_mask;
        fp_bkq_4_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_4_com_2 = 12'h0;
        fp_bkq_4_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_5_com_2;
  wire [11:0] fp_bkq_5_uncom_2;

  always @(*)
  begin
    fp_bkq_5_com_2 = 12'h0;
    fp_bkq_5_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.queue.valids_5 && !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx))
      begin
        fp_bkq_5_com_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_br_mask;
        fp_bkq_5_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_5_com_2 = 12'h0;
        fp_bkq_5_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_6_com_2;
  wire [11:0] fp_bkq_6_uncom_2;

  always @(*)
  begin
    fp_bkq_6_com_2 = 12'h0;
    fp_bkq_6_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.queue.valids_6 && !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx))
      begin
        fp_bkq_6_com_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_br_mask;
        fp_bkq_6_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_6_com_2 = 12'h0;
        fp_bkq_6_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_1_0_com_2;
  wire [11:0] fp_bkq_1_0_uncom_2;

  always @(*)
  begin
    fp_bkq_1_0_com_2 = 12'h0;
    fp_bkq_1_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0 && !(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx))
      begin
        fp_bkq_1_0_com_2 = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_br_mask;
        fp_bkq_1_0_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_1_0_com_2 = 12'h0;
        fp_bkq_1_0_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_1_1_com_2;
  wire [11:0] fp_bkq_1_1_uncom_2;

  always @(*)
  begin
    fp_bkq_1_1_com_2 = 12'h0;
    fp_bkq_1_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1 && !(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx))
      begin
        fp_bkq_1_1_com_2 = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_br_mask;
        fp_bkq_1_1_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_1_1_com_2 = 12'h0;
        fp_bkq_1_1_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_br_mask;
      end
    end
  end

  wire [11:0] fp_bkq_1_2_com_2;
  wire [11:0] fp_bkq_1_2_uncom_2;

  always @(*)
  begin
    fp_bkq_1_2_com_2 = 12'h0;
    fp_bkq_1_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2 && !(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx))
      begin
        fp_bkq_1_2_com_2 = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_br_mask;
        fp_bkq_1_2_uncom_2 = 12'hfff;
      end
      else
      begin
        fp_bkq_1_2_com_2 = 12'h0;
        fp_bkq_1_2_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_br_mask;
      end
    end
  end

  wire [11:0] fdiv_buf_com_2;
  wire [11:0] fdiv_buf_uncom_2;

  always @(*)
  begin
    fdiv_buf_com_2 = 12'h0;
    fdiv_buf_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_val)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx))
      begin
        fdiv_buf_com_2 = soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_br_mask;
        fdiv_buf_uncom_2 = 12'hfff;
      end
      else
      begin
        fdiv_buf_com_2 = 12'h0;
        fdiv_buf_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_br_mask;
      end
    end
  end

  wire [11:0] fdiv_divsqrt_com_2;
  wire [11:0] fdiv_divsqrt_uncom_2;

  always @(*)
  begin
    fdiv_divsqrt_com_2 = 12'h0;
    fdiv_divsqrt_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx))
      begin
        fdiv_divsqrt_com_2 = soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_br_mask;
        fdiv_divsqrt_uncom_2 = 12'hfff;
      end
      else
      begin
        fdiv_divsqrt_com_2 = 12'h0;
        fdiv_divsqrt_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_br_mask;
      end
    end
  end

  wire [11:0] fdiv_out_com_2;
  wire [11:0] fdiv_out_uncom_2;

  always @(*)
  begin
    fdiv_out_com_2 = 12'h0;
    fdiv_out_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_val)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx))
      begin
        fdiv_out_com_2 = soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_br_mask;
        fdiv_out_uncom_2 = 12'hfff;
      end
      else
      begin
        fdiv_out_com_2 = 12'h0;
        fdiv_out_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_br_mask;
      end
    end
  end

  wire [11:0] fpu_T_2_0_com_2;
  wire [11:0] fpu_T_2_0_uncom_2;

  always @(*)
  begin
    fpu_T_2_0_com_2 = 12'h0;
    fpu_T_2_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_0 && !(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx))
      begin
        fpu_T_2_0_com_2 = soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_br_mask;
        fpu_T_2_0_uncom_2 = 12'hfff;
      end
      else
      begin
        fpu_T_2_0_com_2 = 12'h0;
        fpu_T_2_0_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_br_mask;
      end
    end
  end

  wire [11:0] fpu_T_2_1_com_2;
  wire [11:0] fpu_T_2_1_uncom_2;

  always @(*)
  begin
    fpu_T_2_1_com_2 = 12'h0;
    fpu_T_2_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_1 && !(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx))
      begin
        fpu_T_2_1_com_2 = soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_br_mask;
        fpu_T_2_1_uncom_2 = 12'hfff;
      end
      else
      begin
        fpu_T_2_1_com_2 = 12'h0;
        fpu_T_2_1_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_br_mask;
      end
    end
  end

  wire [11:0] fpu_T_2_2_com_2;
  wire [11:0] fpu_T_2_2_uncom_2;

  always @(*)
  begin
    fpu_T_2_2_com_2 = 12'h0;
    fpu_T_2_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_2 && !(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx))
      begin
        fpu_T_2_2_com_2 = soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_br_mask;
        fpu_T_2_2_uncom_2 = 12'hfff;
      end
      else
      begin
        fpu_T_2_2_com_2 = 12'h0;
        fpu_T_2_2_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_br_mask;
      end
    end
  end

  wire [11:0] fpu_T_2_3_com_2;
  wire [11:0] fpu_T_2_3_uncom_2;

  always @(*)
  begin
    fpu_T_2_3_com_2 = 12'h0;
    fpu_T_2_3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx) && soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_3 && !(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx))
      begin
        fpu_T_2_3_com_2 = soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_br_mask;
        fpu_T_2_3_uncom_2 = 12'hfff;
      end
      else
      begin
        fpu_T_2_3_com_2 = 12'h0;
        fpu_T_2_3_uncom_2 = soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_br_mask;
      end
    end
  end

  wire [11:0] f_exe_reg_com_2;
  wire [11:0] f_exe_reg_uncom_2;

  always @(*)
  begin
    f_exe_reg_com_2 = 12'h0;
    f_exe_reg_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx) && soc2.core.fp_pipeline.fregister_read.exe_reg_valids_0 && !(soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx))
      begin
        f_exe_reg_com_2 = soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_br_mask;
        f_exe_reg_uncom_2 = 12'hfff;
      end
      else
      begin
        f_exe_reg_com_2 = 12'h0;
        f_exe_reg_uncom_2 = soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_br_mask;
      end
    end
  end

  wire [11:0] f_rrd_com_2;
  wire [11:0] f_rrd_uncom_2;

  always @(*)
  begin
    f_rrd_com_2 = 12'h0;
    f_rrd_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx) && soc2.core.fp_pipeline.fregister_read.rrd_valids_0_REG && !(soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx))
      begin
        f_rrd_com_2 = soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_br_mask;
        f_rrd_uncom_2 = 12'hfff;
      end
      else
      begin
        f_rrd_com_2 = 12'h0;
        f_rrd_uncom_2 = soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_0_com_2;
  wire [11:0] int_issue_slot_0_uncom_2;

  always @(*)
  begin
    int_issue_slot_0_com_2 = 12'h0;
    int_issue_slot_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_0.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_0.io_valid && !(soc2.core.int_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_0.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_0.slot_uop_rob_idx))
      begin
        int_issue_slot_0_com_2 = soc2.core.int_issue_unit.slots_0.slot_uop_br_mask;
        int_issue_slot_0_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_0_com_2 = 12'h0;
        int_issue_slot_0_uncom_2 = soc2.core.int_issue_unit.slots_0.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_1_com_2;
  wire [11:0] int_issue_slot_1_uncom_2;

  always @(*)
  begin
    int_issue_slot_1_com_2 = 12'h0;
    int_issue_slot_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_1.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_1.io_valid && !(soc2.core.int_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_1.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_1.slot_uop_rob_idx))
      begin
        int_issue_slot_1_com_2 = soc2.core.int_issue_unit.slots_1.slot_uop_br_mask;
        int_issue_slot_1_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_1_com_2 = 12'h0;
        int_issue_slot_1_uncom_2 = soc2.core.int_issue_unit.slots_1.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_2_com_2;
  wire [11:0] int_issue_slot_2_uncom_2;

  always @(*)
  begin
    int_issue_slot_2_com_2 = 12'h0;
    int_issue_slot_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_2.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_2.io_valid && !(soc2.core.int_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_2.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_2.slot_uop_rob_idx))
      begin
        int_issue_slot_2_com_2 = soc2.core.int_issue_unit.slots_2.slot_uop_br_mask;
        int_issue_slot_2_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_2_com_2 = 12'h0;
        int_issue_slot_2_uncom_2 = soc2.core.int_issue_unit.slots_2.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_3_com_2;
  wire [11:0] int_issue_slot_3_uncom_2;

  always @(*)
  begin
    int_issue_slot_3_com_2 = 12'h0;
    int_issue_slot_3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_3.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_3.io_valid && !(soc2.core.int_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_3.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_3.slot_uop_rob_idx))
      begin
        int_issue_slot_3_com_2 = soc2.core.int_issue_unit.slots_3.slot_uop_br_mask;
        int_issue_slot_3_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_3_com_2 = 12'h0;
        int_issue_slot_3_uncom_2 = soc2.core.int_issue_unit.slots_3.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_4_com_2;
  wire [11:0] int_issue_slot_4_uncom_2;

  always @(*)
  begin
    int_issue_slot_4_com_2 = 12'h0;
    int_issue_slot_4_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_4.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_4.io_valid && !(soc2.core.int_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_4.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_4.slot_uop_rob_idx))
      begin
        int_issue_slot_4_com_2 = soc2.core.int_issue_unit.slots_4.slot_uop_br_mask;
        int_issue_slot_4_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_4_com_2 = 12'h0;
        int_issue_slot_4_uncom_2 = soc2.core.int_issue_unit.slots_4.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_5_com_2;
  wire [11:0] int_issue_slot_5_uncom_2;

  always @(*)
  begin
    int_issue_slot_5_com_2 = 12'h0;
    int_issue_slot_5_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_5.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_5.io_valid && !(soc2.core.int_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_5.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_5.slot_uop_rob_idx))
      begin
        int_issue_slot_5_com_2 = soc2.core.int_issue_unit.slots_5.slot_uop_br_mask;
        int_issue_slot_5_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_5_com_2 = 12'h0;
        int_issue_slot_5_uncom_2 = soc2.core.int_issue_unit.slots_5.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_6_com_2;
  wire [11:0] int_issue_slot_6_uncom_2;

  always @(*)
  begin
    int_issue_slot_6_com_2 = 12'h0;
    int_issue_slot_6_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_6.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_6.io_valid && !(soc2.core.int_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_6.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_6.slot_uop_rob_idx))
      begin
        int_issue_slot_6_com_2 = soc2.core.int_issue_unit.slots_6.slot_uop_br_mask;
        int_issue_slot_6_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_6_com_2 = 12'h0;
        int_issue_slot_6_uncom_2 = soc2.core.int_issue_unit.slots_6.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_7_com_2;
  wire [11:0] int_issue_slot_7_uncom_2;

  always @(*)
  begin
    int_issue_slot_7_com_2 = 12'h0;
    int_issue_slot_7_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_7.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_7.io_valid && !(soc2.core.int_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_7.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_7.slot_uop_rob_idx))
      begin
        int_issue_slot_7_com_2 = soc2.core.int_issue_unit.slots_7.slot_uop_br_mask;
        int_issue_slot_7_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_7_com_2 = 12'h0;
        int_issue_slot_7_uncom_2 = soc2.core.int_issue_unit.slots_7.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_8_com_2;
  wire [11:0] int_issue_slot_8_uncom_2;

  always @(*)
  begin
    int_issue_slot_8_com_2 = 12'h0;
    int_issue_slot_8_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_8.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_8.io_valid && !(soc2.core.int_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_8.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_8.slot_uop_rob_idx))
      begin
        int_issue_slot_8_com_2 = soc2.core.int_issue_unit.slots_8.slot_uop_br_mask;
        int_issue_slot_8_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_8_com_2 = 12'h0;
        int_issue_slot_8_uncom_2 = soc2.core.int_issue_unit.slots_8.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_9_com_2;
  wire [11:0] int_issue_slot_9_uncom_2;

  always @(*)
  begin
    int_issue_slot_9_com_2 = 12'h0;
    int_issue_slot_9_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_9.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_9.io_valid && !(soc2.core.int_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_9.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_9.slot_uop_rob_idx))
      begin
        int_issue_slot_9_com_2 = soc2.core.int_issue_unit.slots_9.slot_uop_br_mask;
        int_issue_slot_9_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_9_com_2 = 12'h0;
        int_issue_slot_9_uncom_2 = soc2.core.int_issue_unit.slots_9.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_10_com_2;
  wire [11:0] int_issue_slot_10_uncom_2;

  always @(*)
  begin
    int_issue_slot_10_com_2 = 12'h0;
    int_issue_slot_10_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_10.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_10.io_valid && !(soc2.core.int_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_10.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_10.slot_uop_rob_idx))
      begin
        int_issue_slot_10_com_2 = soc2.core.int_issue_unit.slots_10.slot_uop_br_mask;
        int_issue_slot_10_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_10_com_2 = 12'h0;
        int_issue_slot_10_uncom_2 = soc2.core.int_issue_unit.slots_10.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_11_com_2;
  wire [11:0] int_issue_slot_11_uncom_2;

  always @(*)
  begin
    int_issue_slot_11_com_2 = 12'h0;
    int_issue_slot_11_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_11.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_11.io_valid && !(soc2.core.int_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_11.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_11.slot_uop_rob_idx))
      begin
        int_issue_slot_11_com_2 = soc2.core.int_issue_unit.slots_11.slot_uop_br_mask;
        int_issue_slot_11_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_11_com_2 = 12'h0;
        int_issue_slot_11_uncom_2 = soc2.core.int_issue_unit.slots_11.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_12_com_2;
  wire [11:0] int_issue_slot_12_uncom_2;

  always @(*)
  begin
    int_issue_slot_12_com_2 = 12'h0;
    int_issue_slot_12_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_12.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_12.io_valid && !(soc2.core.int_issue_unit.slots_12.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_12.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_12.slot_uop_rob_idx))
      begin
        int_issue_slot_12_com_2 = soc2.core.int_issue_unit.slots_12.slot_uop_br_mask;
        int_issue_slot_12_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_12_com_2 = 12'h0;
        int_issue_slot_12_uncom_2 = soc2.core.int_issue_unit.slots_12.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_13_com_2;
  wire [11:0] int_issue_slot_13_uncom_2;

  always @(*)
  begin
    int_issue_slot_13_com_2 = 12'h0;
    int_issue_slot_13_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_13.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_13.io_valid && !(soc2.core.int_issue_unit.slots_13.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_13.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_13.slot_uop_rob_idx))
      begin
        int_issue_slot_13_com_2 = soc2.core.int_issue_unit.slots_13.slot_uop_br_mask;
        int_issue_slot_13_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_13_com_2 = 12'h0;
        int_issue_slot_13_uncom_2 = soc2.core.int_issue_unit.slots_13.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_14_com_2;
  wire [11:0] int_issue_slot_14_uncom_2;

  always @(*)
  begin
    int_issue_slot_14_com_2 = 12'h0;
    int_issue_slot_14_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_14.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_14.io_valid && !(soc2.core.int_issue_unit.slots_14.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_14.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_14.slot_uop_rob_idx))
      begin
        int_issue_slot_14_com_2 = soc2.core.int_issue_unit.slots_14.slot_uop_br_mask;
        int_issue_slot_14_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_14_com_2 = 12'h0;
        int_issue_slot_14_uncom_2 = soc2.core.int_issue_unit.slots_14.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_15_com_2;
  wire [11:0] int_issue_slot_15_uncom_2;

  always @(*)
  begin
    int_issue_slot_15_com_2 = 12'h0;
    int_issue_slot_15_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_15.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_15.io_valid && !(soc2.core.int_issue_unit.slots_15.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_15.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_15.slot_uop_rob_idx))
      begin
        int_issue_slot_15_com_2 = soc2.core.int_issue_unit.slots_15.slot_uop_br_mask;
        int_issue_slot_15_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_15_com_2 = 12'h0;
        int_issue_slot_15_uncom_2 = soc2.core.int_issue_unit.slots_15.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_16_com_2;
  wire [11:0] int_issue_slot_16_uncom_2;

  always @(*)
  begin
    int_issue_slot_16_com_2 = 12'h0;
    int_issue_slot_16_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_16.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_16.io_valid && !(soc2.core.int_issue_unit.slots_16.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_16.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_16.slot_uop_rob_idx))
      begin
        int_issue_slot_16_com_2 = soc2.core.int_issue_unit.slots_16.slot_uop_br_mask;
        int_issue_slot_16_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_16_com_2 = 12'h0;
        int_issue_slot_16_uncom_2 = soc2.core.int_issue_unit.slots_16.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_17_com_2;
  wire [11:0] int_issue_slot_17_uncom_2;

  always @(*)
  begin
    int_issue_slot_17_com_2 = 12'h0;
    int_issue_slot_17_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_17.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_17.io_valid && !(soc2.core.int_issue_unit.slots_17.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_17.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_17.slot_uop_rob_idx))
      begin
        int_issue_slot_17_com_2 = soc2.core.int_issue_unit.slots_17.slot_uop_br_mask;
        int_issue_slot_17_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_17_com_2 = 12'h0;
        int_issue_slot_17_uncom_2 = soc2.core.int_issue_unit.slots_17.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_18_com_2;
  wire [11:0] int_issue_slot_18_uncom_2;

  always @(*)
  begin
    int_issue_slot_18_com_2 = 12'h0;
    int_issue_slot_18_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_18.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_18.io_valid && !(soc2.core.int_issue_unit.slots_18.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_18.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_18.slot_uop_rob_idx))
      begin
        int_issue_slot_18_com_2 = soc2.core.int_issue_unit.slots_18.slot_uop_br_mask;
        int_issue_slot_18_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_18_com_2 = 12'h0;
        int_issue_slot_18_uncom_2 = soc2.core.int_issue_unit.slots_18.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] int_issue_slot_19_com_2;
  wire [11:0] int_issue_slot_19_uncom_2;

  always @(*)
  begin
    int_issue_slot_19_com_2 = 12'h0;
    int_issue_slot_19_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.int_issue_unit.slots_19.slot_uop_rob_idx) && soc2.core.int_issue_unit.slots_19.io_valid && !(soc2.core.int_issue_unit.slots_19.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_19.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_19.slot_uop_rob_idx))
      begin
        int_issue_slot_19_com_2 = soc2.core.int_issue_unit.slots_19.slot_uop_br_mask;
        int_issue_slot_19_uncom_2 = 12'hfff;
      end
      else
      begin
        int_issue_slot_19_com_2 = 12'h0;
        int_issue_slot_19_uncom_2 = soc2.core.int_issue_unit.slots_19.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_0_com_2;
  wire [11:0] mem_issue_slot_0_uncom_2;

  always @(*)
  begin
    mem_issue_slot_0_com_2 = 12'h0;
    mem_issue_slot_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_0.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_0.io_valid && !(soc2.core.mem_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_0.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_0.slot_uop_rob_idx))
      begin
        mem_issue_slot_0_com_2 = soc2.core.mem_issue_unit.slots_0.slot_uop_br_mask;
        mem_issue_slot_0_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_0_com_2 = 12'h0;
        mem_issue_slot_0_uncom_2 = soc2.core.mem_issue_unit.slots_0.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_1_com_2;
  wire [11:0] mem_issue_slot_1_uncom_2;

  always @(*)
  begin
    mem_issue_slot_1_com_2 = 12'h0;
    mem_issue_slot_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_1.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_1.io_valid && !(soc2.core.mem_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_1.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_1.slot_uop_rob_idx))
      begin
        mem_issue_slot_1_com_2 = soc2.core.mem_issue_unit.slots_1.slot_uop_br_mask;
        mem_issue_slot_1_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_1_com_2 = 12'h0;
        mem_issue_slot_1_uncom_2 = soc2.core.mem_issue_unit.slots_1.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_2_com_2;
  wire [11:0] mem_issue_slot_2_uncom_2;

  always @(*)
  begin
    mem_issue_slot_2_com_2 = 12'h0;
    mem_issue_slot_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_2.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_2.io_valid && !(soc2.core.mem_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_2.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_2.slot_uop_rob_idx))
      begin
        mem_issue_slot_2_com_2 = soc2.core.mem_issue_unit.slots_2.slot_uop_br_mask;
        mem_issue_slot_2_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_2_com_2 = 12'h0;
        mem_issue_slot_2_uncom_2 = soc2.core.mem_issue_unit.slots_2.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_3_com_2;
  wire [11:0] mem_issue_slot_3_uncom_2;

  always @(*)
  begin
    mem_issue_slot_3_com_2 = 12'h0;
    mem_issue_slot_3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_3.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_3.io_valid && !(soc2.core.mem_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_3.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_3.slot_uop_rob_idx))
      begin
        mem_issue_slot_3_com_2 = soc2.core.mem_issue_unit.slots_3.slot_uop_br_mask;
        mem_issue_slot_3_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_3_com_2 = 12'h0;
        mem_issue_slot_3_uncom_2 = soc2.core.mem_issue_unit.slots_3.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_4_com_2;
  wire [11:0] mem_issue_slot_4_uncom_2;

  always @(*)
  begin
    mem_issue_slot_4_com_2 = 12'h0;
    mem_issue_slot_4_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_4.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_4.io_valid && !(soc2.core.mem_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_4.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_4.slot_uop_rob_idx))
      begin
        mem_issue_slot_4_com_2 = soc2.core.mem_issue_unit.slots_4.slot_uop_br_mask;
        mem_issue_slot_4_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_4_com_2 = 12'h0;
        mem_issue_slot_4_uncom_2 = soc2.core.mem_issue_unit.slots_4.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_5_com_2;
  wire [11:0] mem_issue_slot_5_uncom_2;

  always @(*)
  begin
    mem_issue_slot_5_com_2 = 12'h0;
    mem_issue_slot_5_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_5.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_5.io_valid && !(soc2.core.mem_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_5.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_5.slot_uop_rob_idx))
      begin
        mem_issue_slot_5_com_2 = soc2.core.mem_issue_unit.slots_5.slot_uop_br_mask;
        mem_issue_slot_5_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_5_com_2 = 12'h0;
        mem_issue_slot_5_uncom_2 = soc2.core.mem_issue_unit.slots_5.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_6_com_2;
  wire [11:0] mem_issue_slot_6_uncom_2;

  always @(*)
  begin
    mem_issue_slot_6_com_2 = 12'h0;
    mem_issue_slot_6_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_6.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_6.io_valid && !(soc2.core.mem_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_6.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_6.slot_uop_rob_idx))
      begin
        mem_issue_slot_6_com_2 = soc2.core.mem_issue_unit.slots_6.slot_uop_br_mask;
        mem_issue_slot_6_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_6_com_2 = 12'h0;
        mem_issue_slot_6_uncom_2 = soc2.core.mem_issue_unit.slots_6.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_7_com_2;
  wire [11:0] mem_issue_slot_7_uncom_2;

  always @(*)
  begin
    mem_issue_slot_7_com_2 = 12'h0;
    mem_issue_slot_7_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_7.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_7.io_valid && !(soc2.core.mem_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_7.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_7.slot_uop_rob_idx))
      begin
        mem_issue_slot_7_com_2 = soc2.core.mem_issue_unit.slots_7.slot_uop_br_mask;
        mem_issue_slot_7_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_7_com_2 = 12'h0;
        mem_issue_slot_7_uncom_2 = soc2.core.mem_issue_unit.slots_7.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_8_com_2;
  wire [11:0] mem_issue_slot_8_uncom_2;

  always @(*)
  begin
    mem_issue_slot_8_com_2 = 12'h0;
    mem_issue_slot_8_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_8.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_8.io_valid && !(soc2.core.mem_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_8.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_8.slot_uop_rob_idx))
      begin
        mem_issue_slot_8_com_2 = soc2.core.mem_issue_unit.slots_8.slot_uop_br_mask;
        mem_issue_slot_8_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_8_com_2 = 12'h0;
        mem_issue_slot_8_uncom_2 = soc2.core.mem_issue_unit.slots_8.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_9_com_2;
  wire [11:0] mem_issue_slot_9_uncom_2;

  always @(*)
  begin
    mem_issue_slot_9_com_2 = 12'h0;
    mem_issue_slot_9_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_9.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_9.io_valid && !(soc2.core.mem_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_9.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_9.slot_uop_rob_idx))
      begin
        mem_issue_slot_9_com_2 = soc2.core.mem_issue_unit.slots_9.slot_uop_br_mask;
        mem_issue_slot_9_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_9_com_2 = 12'h0;
        mem_issue_slot_9_uncom_2 = soc2.core.mem_issue_unit.slots_9.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_10_com_2;
  wire [11:0] mem_issue_slot_10_uncom_2;

  always @(*)
  begin
    mem_issue_slot_10_com_2 = 12'h0;
    mem_issue_slot_10_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_10.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_10.io_valid && !(soc2.core.mem_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_10.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_10.slot_uop_rob_idx))
      begin
        mem_issue_slot_10_com_2 = soc2.core.mem_issue_unit.slots_10.slot_uop_br_mask;
        mem_issue_slot_10_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_10_com_2 = 12'h0;
        mem_issue_slot_10_uncom_2 = soc2.core.mem_issue_unit.slots_10.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] mem_issue_slot_11_com_2;
  wire [11:0] mem_issue_slot_11_uncom_2;

  always @(*)
  begin
    mem_issue_slot_11_com_2 = 12'h0;
    mem_issue_slot_11_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.core.mem_issue_unit.slots_11.slot_uop_rob_idx) && soc2.core.mem_issue_unit.slots_11.io_valid && !(soc2.core.mem_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_11.slot_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_11.slot_uop_rob_idx))
      begin
        mem_issue_slot_11_com_2 = soc2.core.mem_issue_unit.slots_11.slot_uop_br_mask;
        mem_issue_slot_11_uncom_2 = 12'hfff;
      end
      else
      begin
        mem_issue_slot_11_com_2 = 12'h0;
        mem_issue_slot_11_uncom_2 = soc2.core.mem_issue_unit.slots_11.slot_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_0_com_2;
  wire [11:0] lsu_ldq_0_uncom_2;

  always @(*)
  begin
    lsu_ldq_0_com_2 = 12'h0;
    lsu_ldq_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_0_bits_uop_rob_idx) && soc2.lsu.ldq_0_valid && !(soc2.lsu.ldq_0_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_0_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_0_bits_uop_rob_idx))
      begin
        lsu_ldq_0_com_2 = soc2.lsu.ldq_0_bits_uop_br_mask;
        lsu_ldq_0_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_0_com_2 = 12'h0;
        lsu_ldq_0_uncom_2 = soc2.lsu.ldq_0_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_1_com_2;
  wire [11:0] lsu_ldq_1_uncom_2;

  always @(*)
  begin
    lsu_ldq_1_com_2 = 12'h0;
    lsu_ldq_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_1_bits_uop_rob_idx) && soc2.lsu.ldq_1_valid && !(soc2.lsu.ldq_1_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_1_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_1_bits_uop_rob_idx))
      begin
        lsu_ldq_1_com_2 = soc2.lsu.ldq_1_bits_uop_br_mask;
        lsu_ldq_1_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_1_com_2 = 12'h0;
        lsu_ldq_1_uncom_2 = soc2.lsu.ldq_1_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_2_com_2;
  wire [11:0] lsu_ldq_2_uncom_2;

  always @(*)
  begin
    lsu_ldq_2_com_2 = 12'h0;
    lsu_ldq_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_2_bits_uop_rob_idx) && soc2.lsu.ldq_2_valid && !(soc2.lsu.ldq_2_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_2_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_2_bits_uop_rob_idx))
      begin
        lsu_ldq_2_com_2 = soc2.lsu.ldq_2_bits_uop_br_mask;
        lsu_ldq_2_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_2_com_2 = 12'h0;
        lsu_ldq_2_uncom_2 = soc2.lsu.ldq_2_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_3_com_2;
  wire [11:0] lsu_ldq_3_uncom_2;

  always @(*)
  begin
    lsu_ldq_3_com_2 = 12'h0;
    lsu_ldq_3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_3_bits_uop_rob_idx) && soc2.lsu.ldq_3_valid && !(soc2.lsu.ldq_3_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_3_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_3_bits_uop_rob_idx))
      begin
        lsu_ldq_3_com_2 = soc2.lsu.ldq_3_bits_uop_br_mask;
        lsu_ldq_3_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_3_com_2 = 12'h0;
        lsu_ldq_3_uncom_2 = soc2.lsu.ldq_3_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_4_com_2;
  wire [11:0] lsu_ldq_4_uncom_2;

  always @(*)
  begin
    lsu_ldq_4_com_2 = 12'h0;
    lsu_ldq_4_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_4_bits_uop_rob_idx) && soc2.lsu.ldq_4_valid && !(soc2.lsu.ldq_4_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_4_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_4_bits_uop_rob_idx))
      begin
        lsu_ldq_4_com_2 = soc2.lsu.ldq_4_bits_uop_br_mask;
        lsu_ldq_4_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_4_com_2 = 12'h0;
        lsu_ldq_4_uncom_2 = soc2.lsu.ldq_4_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_5_com_2;
  wire [11:0] lsu_ldq_5_uncom_2;

  always @(*)
  begin
    lsu_ldq_5_com_2 = 12'h0;
    lsu_ldq_5_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_5_bits_uop_rob_idx) && soc2.lsu.ldq_5_valid && !(soc2.lsu.ldq_5_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_5_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_5_bits_uop_rob_idx))
      begin
        lsu_ldq_5_com_2 = soc2.lsu.ldq_5_bits_uop_br_mask;
        lsu_ldq_5_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_5_com_2 = 12'h0;
        lsu_ldq_5_uncom_2 = soc2.lsu.ldq_5_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_6_com_2;
  wire [11:0] lsu_ldq_6_uncom_2;

  always @(*)
  begin
    lsu_ldq_6_com_2 = 12'h0;
    lsu_ldq_6_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_6_bits_uop_rob_idx) && soc2.lsu.ldq_6_valid && !(soc2.lsu.ldq_6_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_6_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_6_bits_uop_rob_idx))
      begin
        lsu_ldq_6_com_2 = soc2.lsu.ldq_6_bits_uop_br_mask;
        lsu_ldq_6_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_6_com_2 = 12'h0;
        lsu_ldq_6_uncom_2 = soc2.lsu.ldq_6_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_7_com_2;
  wire [11:0] lsu_ldq_7_uncom_2;

  always @(*)
  begin
    lsu_ldq_7_com_2 = 12'h0;
    lsu_ldq_7_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_7_bits_uop_rob_idx) && soc2.lsu.ldq_7_valid && !(soc2.lsu.ldq_7_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_7_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_7_bits_uop_rob_idx))
      begin
        lsu_ldq_7_com_2 = soc2.lsu.ldq_7_bits_uop_br_mask;
        lsu_ldq_7_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_7_com_2 = 12'h0;
        lsu_ldq_7_uncom_2 = soc2.lsu.ldq_7_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_8_com_2;
  wire [11:0] lsu_ldq_8_uncom_2;

  always @(*)
  begin
    lsu_ldq_8_com_2 = 12'h0;
    lsu_ldq_8_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_8_bits_uop_rob_idx) && soc2.lsu.ldq_8_valid && !(soc2.lsu.ldq_8_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_8_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_8_bits_uop_rob_idx))
      begin
        lsu_ldq_8_com_2 = soc2.lsu.ldq_8_bits_uop_br_mask;
        lsu_ldq_8_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_8_com_2 = 12'h0;
        lsu_ldq_8_uncom_2 = soc2.lsu.ldq_8_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_9_com_2;
  wire [11:0] lsu_ldq_9_uncom_2;

  always @(*)
  begin
    lsu_ldq_9_com_2 = 12'h0;
    lsu_ldq_9_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_9_bits_uop_rob_idx) && soc2.lsu.ldq_9_valid && !(soc2.lsu.ldq_9_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_9_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_9_bits_uop_rob_idx))
      begin
        lsu_ldq_9_com_2 = soc2.lsu.ldq_9_bits_uop_br_mask;
        lsu_ldq_9_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_9_com_2 = 12'h0;
        lsu_ldq_9_uncom_2 = soc2.lsu.ldq_9_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_10_com_2;
  wire [11:0] lsu_ldq_10_uncom_2;

  always @(*)
  begin
    lsu_ldq_10_com_2 = 12'h0;
    lsu_ldq_10_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_10_bits_uop_rob_idx) && soc2.lsu.ldq_10_valid && !(soc2.lsu.ldq_10_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_10_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_10_bits_uop_rob_idx))
      begin
        lsu_ldq_10_com_2 = soc2.lsu.ldq_10_bits_uop_br_mask;
        lsu_ldq_10_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_10_com_2 = 12'h0;
        lsu_ldq_10_uncom_2 = soc2.lsu.ldq_10_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_11_com_2;
  wire [11:0] lsu_ldq_11_uncom_2;

  always @(*)
  begin
    lsu_ldq_11_com_2 = 12'h0;
    lsu_ldq_11_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_11_bits_uop_rob_idx) && soc2.lsu.ldq_11_valid && !(soc2.lsu.ldq_11_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_11_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_11_bits_uop_rob_idx))
      begin
        lsu_ldq_11_com_2 = soc2.lsu.ldq_11_bits_uop_br_mask;
        lsu_ldq_11_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_11_com_2 = 12'h0;
        lsu_ldq_11_uncom_2 = soc2.lsu.ldq_11_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_12_com_2;
  wire [11:0] lsu_ldq_12_uncom_2;

  always @(*)
  begin
    lsu_ldq_12_com_2 = 12'h0;
    lsu_ldq_12_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_12_bits_uop_rob_idx) && soc2.lsu.ldq_12_valid && !(soc2.lsu.ldq_12_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_12_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_12_bits_uop_rob_idx))
      begin
        lsu_ldq_12_com_2 = soc2.lsu.ldq_12_bits_uop_br_mask;
        lsu_ldq_12_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_12_com_2 = 12'h0;
        lsu_ldq_12_uncom_2 = soc2.lsu.ldq_12_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_13_com_2;
  wire [11:0] lsu_ldq_13_uncom_2;

  always @(*)
  begin
    lsu_ldq_13_com_2 = 12'h0;
    lsu_ldq_13_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_13_bits_uop_rob_idx) && soc2.lsu.ldq_13_valid && !(soc2.lsu.ldq_13_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_13_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_13_bits_uop_rob_idx))
      begin
        lsu_ldq_13_com_2 = soc2.lsu.ldq_13_bits_uop_br_mask;
        lsu_ldq_13_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_13_com_2 = 12'h0;
        lsu_ldq_13_uncom_2 = soc2.lsu.ldq_13_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_14_com_2;
  wire [11:0] lsu_ldq_14_uncom_2;

  always @(*)
  begin
    lsu_ldq_14_com_2 = 12'h0;
    lsu_ldq_14_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_14_bits_uop_rob_idx) && soc2.lsu.ldq_14_valid && !(soc2.lsu.ldq_14_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_14_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_14_bits_uop_rob_idx))
      begin
        lsu_ldq_14_com_2 = soc2.lsu.ldq_14_bits_uop_br_mask;
        lsu_ldq_14_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_14_com_2 = 12'h0;
        lsu_ldq_14_uncom_2 = soc2.lsu.ldq_14_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_ldq_15_com_2;
  wire [11:0] lsu_ldq_15_uncom_2;

  always @(*)
  begin
    lsu_ldq_15_com_2 = 12'h0;
    lsu_ldq_15_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.ldq_15_bits_uop_rob_idx) && soc2.lsu.ldq_15_valid && !(soc2.lsu.ldq_15_bits_uop_uses_stq && stq_committed_2[soc2.lsu.ldq_15_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_15_bits_uop_rob_idx))
      begin
        lsu_ldq_15_com_2 = soc2.lsu.ldq_15_bits_uop_br_mask;
        lsu_ldq_15_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_ldq_15_com_2 = 12'h0;
        lsu_ldq_15_uncom_2 = soc2.lsu.ldq_15_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_com_2;
  wire [11:0] lsu_mem_uncom_2;

  always @(*)
  begin
    lsu_mem_com_2 = 12'h0;
    lsu_mem_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.mem_incoming_uop_0_rob_idx) && soc2.lsu.fired_sfence_0)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.mem_incoming_uop_0_rob_idx))
      begin
        lsu_mem_com_2 = soc2.lsu.mem_incoming_uop_0_br_mask;
        lsu_mem_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_mem_com_2 = 12'h0;
        lsu_mem_uncom_2 = soc2.lsu.mem_incoming_uop_0_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_stq_com_2;
  wire [11:0] lsu_mem_stq_uncom_2;

  always @(*)
  begin
    lsu_mem_stq_com_2 = 12'h0;
    lsu_mem_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx) && (soc2.lsu.fired_stad_incoming_REG || soc2.lsu.fired_sta_incoming_REG || soc2.lsu.fired_std_incoming_REG) && !(stq_committed_2[soc2.lsu.mem_stq_incoming_e_0_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx))
      begin
        lsu_mem_stq_com_2 = soc2.lsu.mem_stq_incoming_e_0_bits_uop_br_mask;
        lsu_mem_stq_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_mem_stq_com_2 = 12'h0;
        lsu_mem_stq_uncom_2 = soc2.lsu.mem_stq_incoming_e_0_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_retry_com_2;
  wire [11:0] lsu_mem_retry_uncom_2;

  always @(*)
  begin
    lsu_mem_retry_com_2 = 12'h0;
    lsu_mem_retry_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.mem_stq_retry_e_bits_uop_rob_idx) && soc2.lsu.fired_sta_retry_REG && !(stq_committed_2[soc2.lsu.mem_stq_retry_e_bits_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.mem_stq_retry_e_bits_uop_rob_idx))
      begin
        lsu_mem_retry_com_2 = soc2.lsu.mem_stq_retry_e_bits_uop_br_mask;
        lsu_mem_retry_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_mem_retry_com_2 = 12'h0;
        lsu_mem_retry_uncom_2 = soc2.lsu.mem_stq_retry_e_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_xcpt_com_2;
  wire [11:0] lsu_mem_xcpt_uncom_2;

  always @(*)
  begin
    lsu_mem_xcpt_com_2 = 12'h0;
    lsu_mem_xcpt_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.mem_xcpt_uops_0_rob_idx) && soc2.lsu.mem_xcpt_valids_0 && !(soc2.lsu.mem_xcpt_uops_0_uses_stq && stq_committed_2[soc2.lsu.mem_xcpt_uops_0_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.mem_xcpt_uops_0_rob_idx))
      begin
        lsu_mem_xcpt_com_2 = soc2.lsu.mem_xcpt_uops_0_br_mask;
        lsu_mem_xcpt_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_mem_xcpt_com_2 = 12'h0;
        lsu_mem_xcpt_uncom_2 = soc2.lsu.mem_xcpt_uops_0_br_mask;
      end
    end
  end

  wire [11:0] lsu_mem_stdf_com_2;
  wire [11:0] lsu_mem_stdf_uncom_2;

  always @(*)
  begin
    lsu_mem_stdf_com_2 = 12'h0;
    lsu_mem_stdf_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.mem_stdf_uop_rob_idx) && soc2.lsu.fired_stdf_incoming && !(stq_committed_2[soc2.lsu.mem_stdf_uop_stq_idx]))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.mem_stdf_uop_rob_idx))
      begin
        lsu_mem_stdf_com_2 = soc2.lsu.mem_stdf_uop_br_mask;
        lsu_mem_stdf_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_mem_stdf_com_2 = 12'h0;
        lsu_mem_stdf_uncom_2 = soc2.lsu.mem_stdf_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stdf_com_2;
  wire [11:0] lsu_stdf_uncom_2;

  always @(*)
  begin
    lsu_stdf_com_2 = 12'h0;
    lsu_stdf_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stdf_clr_bsy_rob_idx) && soc2.lsu.stdf_clr_bsy_valid)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stdf_clr_bsy_rob_idx))
      begin
        lsu_stdf_com_2 = soc2.lsu.stdf_clr_bsy_brmask;
        lsu_stdf_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stdf_com_2 = 12'h0;
        lsu_stdf_uncom_2 = soc2.lsu.stdf_clr_bsy_brmask;
      end
    end
  end

  wire [11:0] lsu_stq_0_com_2;
  wire [11:0] lsu_stq_0_uncom_2;

  always @(*)
  begin
    lsu_stq_0_com_2 = 12'h0;
    lsu_stq_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_0_bits_uop_rob_idx) && soc2.lsu.stq_0_valid && !soc2.lsu.stq_0_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_0_bits_uop_rob_idx))
      begin
        lsu_stq_0_com_2 = soc2.lsu.stq_0_bits_uop_br_mask;
        lsu_stq_0_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_0_com_2 = 12'h0;
        lsu_stq_0_uncom_2 = soc2.lsu.stq_0_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_1_com_2;
  wire [11:0] lsu_stq_1_uncom_2;

  always @(*)
  begin
    lsu_stq_1_com_2 = 12'h0;
    lsu_stq_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_1_bits_uop_rob_idx) && soc2.lsu.stq_1_valid && !soc2.lsu.stq_1_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_1_bits_uop_rob_idx))
      begin
        lsu_stq_1_com_2 = soc2.lsu.stq_1_bits_uop_br_mask;
        lsu_stq_1_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_1_com_2 = 12'h0;
        lsu_stq_1_uncom_2 = soc2.lsu.stq_1_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_2_com_2;
  wire [11:0] lsu_stq_2_uncom_2;

  always @(*)
  begin
    lsu_stq_2_com_2 = 12'h0;
    lsu_stq_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_2_bits_uop_rob_idx) && soc2.lsu.stq_2_valid && !soc2.lsu.stq_2_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_2_bits_uop_rob_idx))
      begin
        lsu_stq_2_com_2 = soc2.lsu.stq_2_bits_uop_br_mask;
        lsu_stq_2_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_2_com_2 = 12'h0;
        lsu_stq_2_uncom_2 = soc2.lsu.stq_2_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_3_com_2;
  wire [11:0] lsu_stq_3_uncom_2;

  always @(*)
  begin
    lsu_stq_3_com_2 = 12'h0;
    lsu_stq_3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_3_bits_uop_rob_idx) && soc2.lsu.stq_3_valid && !soc2.lsu.stq_3_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_3_bits_uop_rob_idx))
      begin
        lsu_stq_3_com_2 = soc2.lsu.stq_3_bits_uop_br_mask;
        lsu_stq_3_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_3_com_2 = 12'h0;
        lsu_stq_3_uncom_2 = soc2.lsu.stq_3_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_4_com_2;
  wire [11:0] lsu_stq_4_uncom_2;

  always @(*)
  begin
    lsu_stq_4_com_2 = 12'h0;
    lsu_stq_4_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_4_bits_uop_rob_idx) && soc2.lsu.stq_4_valid && !soc2.lsu.stq_4_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_4_bits_uop_rob_idx))
      begin
        lsu_stq_4_com_2 = soc2.lsu.stq_4_bits_uop_br_mask;
        lsu_stq_4_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_4_com_2 = 12'h0;
        lsu_stq_4_uncom_2 = soc2.lsu.stq_4_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_5_com_2;
  wire [11:0] lsu_stq_5_uncom_2;

  always @(*)
  begin
    lsu_stq_5_com_2 = 12'h0;
    lsu_stq_5_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_5_bits_uop_rob_idx) && soc2.lsu.stq_5_valid && !soc2.lsu.stq_5_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_5_bits_uop_rob_idx))
      begin
        lsu_stq_5_com_2 = soc2.lsu.stq_5_bits_uop_br_mask;
        lsu_stq_5_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_5_com_2 = 12'h0;
        lsu_stq_5_uncom_2 = soc2.lsu.stq_5_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_6_com_2;
  wire [11:0] lsu_stq_6_uncom_2;

  always @(*)
  begin
    lsu_stq_6_com_2 = 12'h0;
    lsu_stq_6_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_6_bits_uop_rob_idx) && soc2.lsu.stq_6_valid && !soc2.lsu.stq_6_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_6_bits_uop_rob_idx))
      begin
        lsu_stq_6_com_2 = soc2.lsu.stq_6_bits_uop_br_mask;
        lsu_stq_6_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_6_com_2 = 12'h0;
        lsu_stq_6_uncom_2 = soc2.lsu.stq_6_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_7_com_2;
  wire [11:0] lsu_stq_7_uncom_2;

  always @(*)
  begin
    lsu_stq_7_com_2 = 12'h0;
    lsu_stq_7_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_7_bits_uop_rob_idx) && soc2.lsu.stq_7_valid && !soc2.lsu.stq_7_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_7_bits_uop_rob_idx))
      begin
        lsu_stq_7_com_2 = soc2.lsu.stq_7_bits_uop_br_mask;
        lsu_stq_7_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_7_com_2 = 12'h0;
        lsu_stq_7_uncom_2 = soc2.lsu.stq_7_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_8_com_2;
  wire [11:0] lsu_stq_8_uncom_2;

  always @(*)
  begin
    lsu_stq_8_com_2 = 12'h0;
    lsu_stq_8_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_8_bits_uop_rob_idx) && soc2.lsu.stq_8_valid && !soc2.lsu.stq_8_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_8_bits_uop_rob_idx))
      begin
        lsu_stq_8_com_2 = soc2.lsu.stq_8_bits_uop_br_mask;
        lsu_stq_8_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_8_com_2 = 12'h0;
        lsu_stq_8_uncom_2 = soc2.lsu.stq_8_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_9_com_2;
  wire [11:0] lsu_stq_9_uncom_2;

  always @(*)
  begin
    lsu_stq_9_com_2 = 12'h0;
    lsu_stq_9_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_9_bits_uop_rob_idx) && soc2.lsu.stq_9_valid && !soc2.lsu.stq_9_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_9_bits_uop_rob_idx))
      begin
        lsu_stq_9_com_2 = soc2.lsu.stq_9_bits_uop_br_mask;
        lsu_stq_9_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_9_com_2 = 12'h0;
        lsu_stq_9_uncom_2 = soc2.lsu.stq_9_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_10_com_2;
  wire [11:0] lsu_stq_10_uncom_2;

  always @(*)
  begin
    lsu_stq_10_com_2 = 12'h0;
    lsu_stq_10_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_10_bits_uop_rob_idx) && soc2.lsu.stq_10_valid && !soc2.lsu.stq_10_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_10_bits_uop_rob_idx))
      begin
        lsu_stq_10_com_2 = soc2.lsu.stq_10_bits_uop_br_mask;
        lsu_stq_10_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_10_com_2 = 12'h0;
        lsu_stq_10_uncom_2 = soc2.lsu.stq_10_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_11_com_2;
  wire [11:0] lsu_stq_11_uncom_2;

  always @(*)
  begin
    lsu_stq_11_com_2 = 12'h0;
    lsu_stq_11_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_11_bits_uop_rob_idx) && soc2.lsu.stq_11_valid && !soc2.lsu.stq_11_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_11_bits_uop_rob_idx))
      begin
        lsu_stq_11_com_2 = soc2.lsu.stq_11_bits_uop_br_mask;
        lsu_stq_11_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_11_com_2 = 12'h0;
        lsu_stq_11_uncom_2 = soc2.lsu.stq_11_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_12_com_2;
  wire [11:0] lsu_stq_12_uncom_2;

  always @(*)
  begin
    lsu_stq_12_com_2 = 12'h0;
    lsu_stq_12_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_12_bits_uop_rob_idx) && soc2.lsu.stq_12_valid && !soc2.lsu.stq_12_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_12_bits_uop_rob_idx))
      begin
        lsu_stq_12_com_2 = soc2.lsu.stq_12_bits_uop_br_mask;
        lsu_stq_12_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_12_com_2 = 12'h0;
        lsu_stq_12_uncom_2 = soc2.lsu.stq_12_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_13_com_2;
  wire [11:0] lsu_stq_13_uncom_2;

  always @(*)
  begin
    lsu_stq_13_com_2 = 12'h0;
    lsu_stq_13_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_13_bits_uop_rob_idx) && soc2.lsu.stq_13_valid && !soc2.lsu.stq_13_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_13_bits_uop_rob_idx))
      begin
        lsu_stq_13_com_2 = soc2.lsu.stq_13_bits_uop_br_mask;
        lsu_stq_13_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_13_com_2 = 12'h0;
        lsu_stq_13_uncom_2 = soc2.lsu.stq_13_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_14_com_2;
  wire [11:0] lsu_stq_14_uncom_2;

  always @(*)
  begin
    lsu_stq_14_com_2 = 12'h0;
    lsu_stq_14_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_14_bits_uop_rob_idx) && soc2.lsu.stq_14_valid && !soc2.lsu.stq_14_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_14_bits_uop_rob_idx))
      begin
        lsu_stq_14_com_2 = soc2.lsu.stq_14_bits_uop_br_mask;
        lsu_stq_14_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_14_com_2 = 12'h0;
        lsu_stq_14_uncom_2 = soc2.lsu.stq_14_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] lsu_stq_15_com_2;
  wire [11:0] lsu_stq_15_uncom_2;

  always @(*)
  begin
    lsu_stq_15_com_2 = 12'h0;
    lsu_stq_15_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.stq_15_bits_uop_rob_idx) && soc2.lsu.stq_15_valid && !soc2.lsu.stq_15_bits_committed)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_15_bits_uop_rob_idx))
      begin
        lsu_stq_15_com_2 = soc2.lsu.stq_15_bits_uop_br_mask;
        lsu_stq_15_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_stq_15_com_2 = 12'h0;
        lsu_stq_15_uncom_2 = soc2.lsu.stq_15_bits_uop_br_mask;
      end
    end
  end

  wire [11:0] rob__0_com_2;
  wire [11:0] rob__0_uncom_2;

  always @(*)
  begin
    rob__0_com_2 = 12'h0;
    rob__0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b000000))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000000))
      begin
        rob__0_com_2 = soc2.core.rob.rob_uop__0_br_mask;
        rob__0_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__0_com_2 = 12'h0;
        rob__0_uncom_2 = soc2.core.rob.rob_uop__0_br_mask;
      end
    end
  end

  wire [11:0] rob__1_com_2;
  wire [11:0] rob__1_uncom_2;

  always @(*)
  begin
    rob__1_com_2 = 12'h0;
    rob__1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b000010))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000010))
      begin
        rob__1_com_2 = soc2.core.rob.rob_uop__1_br_mask;
        rob__1_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__1_com_2 = 12'h0;
        rob__1_uncom_2 = soc2.core.rob.rob_uop__1_br_mask;
      end
    end
  end

  wire [11:0] rob__2_com_2;
  wire [11:0] rob__2_uncom_2;

  always @(*)
  begin
    rob__2_com_2 = 12'h0;
    rob__2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b000100))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000100))
      begin
        rob__2_com_2 = soc2.core.rob.rob_uop__2_br_mask;
        rob__2_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__2_com_2 = 12'h0;
        rob__2_uncom_2 = soc2.core.rob.rob_uop__2_br_mask;
      end
    end
  end

  wire [11:0] rob__3_com_2;
  wire [11:0] rob__3_uncom_2;

  always @(*)
  begin
    rob__3_com_2 = 12'h0;
    rob__3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b000110))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000110))
      begin
        rob__3_com_2 = soc2.core.rob.rob_uop__3_br_mask;
        rob__3_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__3_com_2 = 12'h0;
        rob__3_uncom_2 = soc2.core.rob.rob_uop__3_br_mask;
      end
    end
  end

  wire [11:0] rob__4_com_2;
  wire [11:0] rob__4_uncom_2;

  always @(*)
  begin
    rob__4_com_2 = 12'h0;
    rob__4_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b001000))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001000))
      begin
        rob__4_com_2 = soc2.core.rob.rob_uop__4_br_mask;
        rob__4_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__4_com_2 = 12'h0;
        rob__4_uncom_2 = soc2.core.rob.rob_uop__4_br_mask;
      end
    end
  end

  wire [11:0] rob__5_com_2;
  wire [11:0] rob__5_uncom_2;

  always @(*)
  begin
    rob__5_com_2 = 12'h0;
    rob__5_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b001010))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001010))
      begin
        rob__5_com_2 = soc2.core.rob.rob_uop__5_br_mask;
        rob__5_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__5_com_2 = 12'h0;
        rob__5_uncom_2 = soc2.core.rob.rob_uop__5_br_mask;
      end
    end
  end

  wire [11:0] rob__6_com_2;
  wire [11:0] rob__6_uncom_2;

  always @(*)
  begin
    rob__6_com_2 = 12'h0;
    rob__6_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b001100))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001100))
      begin
        rob__6_com_2 = soc2.core.rob.rob_uop__6_br_mask;
        rob__6_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__6_com_2 = 12'h0;
        rob__6_uncom_2 = soc2.core.rob.rob_uop__6_br_mask;
      end
    end
  end

  wire [11:0] rob__7_com_2;
  wire [11:0] rob__7_uncom_2;

  always @(*)
  begin
    rob__7_com_2 = 12'h0;
    rob__7_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b001110))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001110))
      begin
        rob__7_com_2 = soc2.core.rob.rob_uop__7_br_mask;
        rob__7_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__7_com_2 = 12'h0;
        rob__7_uncom_2 = soc2.core.rob.rob_uop__7_br_mask;
      end
    end
  end

  wire [11:0] rob__8_com_2;
  wire [11:0] rob__8_uncom_2;

  always @(*)
  begin
    rob__8_com_2 = 12'h0;
    rob__8_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b010000))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010000))
      begin
        rob__8_com_2 = soc2.core.rob.rob_uop__8_br_mask;
        rob__8_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__8_com_2 = 12'h0;
        rob__8_uncom_2 = soc2.core.rob.rob_uop__8_br_mask;
      end
    end
  end

  wire [11:0] rob__9_com_2;
  wire [11:0] rob__9_uncom_2;

  always @(*)
  begin
    rob__9_com_2 = 12'h0;
    rob__9_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b010010))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010010))
      begin
        rob__9_com_2 = soc2.core.rob.rob_uop__9_br_mask;
        rob__9_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__9_com_2 = 12'h0;
        rob__9_uncom_2 = soc2.core.rob.rob_uop__9_br_mask;
      end
    end
  end

  wire [11:0] rob__10_com_2;
  wire [11:0] rob__10_uncom_2;

  always @(*)
  begin
    rob__10_com_2 = 12'h0;
    rob__10_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b010100))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010100))
      begin
        rob__10_com_2 = soc2.core.rob.rob_uop__10_br_mask;
        rob__10_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__10_com_2 = 12'h0;
        rob__10_uncom_2 = soc2.core.rob.rob_uop__10_br_mask;
      end
    end
  end

  wire [11:0] rob__11_com_2;
  wire [11:0] rob__11_uncom_2;

  always @(*)
  begin
    rob__11_com_2 = 12'h0;
    rob__11_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b010110))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010110))
      begin
        rob__11_com_2 = soc2.core.rob.rob_uop__11_br_mask;
        rob__11_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__11_com_2 = 12'h0;
        rob__11_uncom_2 = soc2.core.rob.rob_uop__11_br_mask;
      end
    end
  end

  wire [11:0] rob__12_com_2;
  wire [11:0] rob__12_uncom_2;

  always @(*)
  begin
    rob__12_com_2 = 12'h0;
    rob__12_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b011000))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011000))
      begin
        rob__12_com_2 = soc2.core.rob.rob_uop__12_br_mask;
        rob__12_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__12_com_2 = 12'h0;
        rob__12_uncom_2 = soc2.core.rob.rob_uop__12_br_mask;
      end
    end
  end

  wire [11:0] rob__13_com_2;
  wire [11:0] rob__13_uncom_2;

  always @(*)
  begin
    rob__13_com_2 = 12'h0;
    rob__13_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b011010))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011010))
      begin
        rob__13_com_2 = soc2.core.rob.rob_uop__13_br_mask;
        rob__13_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__13_com_2 = 12'h0;
        rob__13_uncom_2 = soc2.core.rob.rob_uop__13_br_mask;
      end
    end
  end

  wire [11:0] rob__14_com_2;
  wire [11:0] rob__14_uncom_2;

  always @(*)
  begin
    rob__14_com_2 = 12'h0;
    rob__14_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b011100))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011100))
      begin
        rob__14_com_2 = soc2.core.rob.rob_uop__14_br_mask;
        rob__14_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__14_com_2 = 12'h0;
        rob__14_uncom_2 = soc2.core.rob.rob_uop__14_br_mask;
      end
    end
  end

  wire [11:0] rob__15_com_2;
  wire [11:0] rob__15_uncom_2;

  always @(*)
  begin
    rob__15_com_2 = 12'h0;
    rob__15_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b011110))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011110))
      begin
        rob__15_com_2 = soc2.core.rob.rob_uop__15_br_mask;
        rob__15_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__15_com_2 = 12'h0;
        rob__15_uncom_2 = soc2.core.rob.rob_uop__15_br_mask;
      end
    end
  end

  wire [11:0] rob__16_com_2;
  wire [11:0] rob__16_uncom_2;

  always @(*)
  begin
    rob__16_com_2 = 12'h0;
    rob__16_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b100000))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100000))
      begin
        rob__16_com_2 = soc2.core.rob.rob_uop__16_br_mask;
        rob__16_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__16_com_2 = 12'h0;
        rob__16_uncom_2 = soc2.core.rob.rob_uop__16_br_mask;
      end
    end
  end

  wire [11:0] rob__17_com_2;
  wire [11:0] rob__17_uncom_2;

  always @(*)
  begin
    rob__17_com_2 = 12'h0;
    rob__17_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b100010))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100010))
      begin
        rob__17_com_2 = soc2.core.rob.rob_uop__17_br_mask;
        rob__17_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__17_com_2 = 12'h0;
        rob__17_uncom_2 = soc2.core.rob.rob_uop__17_br_mask;
      end
    end
  end

  wire [11:0] rob__18_com_2;
  wire [11:0] rob__18_uncom_2;

  always @(*)
  begin
    rob__18_com_2 = 12'h0;
    rob__18_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b100100))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100100))
      begin
        rob__18_com_2 = soc2.core.rob.rob_uop__18_br_mask;
        rob__18_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__18_com_2 = 12'h0;
        rob__18_uncom_2 = soc2.core.rob.rob_uop__18_br_mask;
      end
    end
  end

  wire [11:0] rob__19_com_2;
  wire [11:0] rob__19_uncom_2;

  always @(*)
  begin
    rob__19_com_2 = 12'h0;
    rob__19_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b100110))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100110))
      begin
        rob__19_com_2 = soc2.core.rob.rob_uop__19_br_mask;
        rob__19_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__19_com_2 = 12'h0;
        rob__19_uncom_2 = soc2.core.rob.rob_uop__19_br_mask;
      end
    end
  end

  wire [11:0] rob__20_com_2;
  wire [11:0] rob__20_uncom_2;

  always @(*)
  begin
    rob__20_com_2 = 12'h0;
    rob__20_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b101000))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101000))
      begin
        rob__20_com_2 = soc2.core.rob.rob_uop__20_br_mask;
        rob__20_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__20_com_2 = 12'h0;
        rob__20_uncom_2 = soc2.core.rob.rob_uop__20_br_mask;
      end
    end
  end

  wire [11:0] rob__21_com_2;
  wire [11:0] rob__21_uncom_2;

  always @(*)
  begin
    rob__21_com_2 = 12'h0;
    rob__21_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b101010))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101010))
      begin
        rob__21_com_2 = soc2.core.rob.rob_uop__21_br_mask;
        rob__21_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__21_com_2 = 12'h0;
        rob__21_uncom_2 = soc2.core.rob.rob_uop__21_br_mask;
      end
    end
  end

  wire [11:0] rob__22_com_2;
  wire [11:0] rob__22_uncom_2;

  always @(*)
  begin
    rob__22_com_2 = 12'h0;
    rob__22_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b101100))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101100))
      begin
        rob__22_com_2 = soc2.core.rob.rob_uop__22_br_mask;
        rob__22_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__22_com_2 = 12'h0;
        rob__22_uncom_2 = soc2.core.rob.rob_uop__22_br_mask;
      end
    end
  end

  wire [11:0] rob__23_com_2;
  wire [11:0] rob__23_uncom_2;

  always @(*)
  begin
    rob__23_com_2 = 12'h0;
    rob__23_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b101110))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101110))
      begin
        rob__23_com_2 = soc2.core.rob.rob_uop__23_br_mask;
        rob__23_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__23_com_2 = 12'h0;
        rob__23_uncom_2 = soc2.core.rob.rob_uop__23_br_mask;
      end
    end
  end

  wire [11:0] rob__24_com_2;
  wire [11:0] rob__24_uncom_2;

  always @(*)
  begin
    rob__24_com_2 = 12'h0;
    rob__24_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b110000))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110000))
      begin
        rob__24_com_2 = soc2.core.rob.rob_uop__24_br_mask;
        rob__24_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__24_com_2 = 12'h0;
        rob__24_uncom_2 = soc2.core.rob.rob_uop__24_br_mask;
      end
    end
  end

  wire [11:0] rob__25_com_2;
  wire [11:0] rob__25_uncom_2;

  always @(*)
  begin
    rob__25_com_2 = 12'h0;
    rob__25_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b110010))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110010))
      begin
        rob__25_com_2 = soc2.core.rob.rob_uop__25_br_mask;
        rob__25_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__25_com_2 = 12'h0;
        rob__25_uncom_2 = soc2.core.rob.rob_uop__25_br_mask;
      end
    end
  end

  wire [11:0] rob__26_com_2;
  wire [11:0] rob__26_uncom_2;

  always @(*)
  begin
    rob__26_com_2 = 12'h0;
    rob__26_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b110100))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110100))
      begin
        rob__26_com_2 = soc2.core.rob.rob_uop__26_br_mask;
        rob__26_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__26_com_2 = 12'h0;
        rob__26_uncom_2 = soc2.core.rob.rob_uop__26_br_mask;
      end
    end
  end

  wire [11:0] rob__27_com_2;
  wire [11:0] rob__27_uncom_2;

  always @(*)
  begin
    rob__27_com_2 = 12'h0;
    rob__27_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b110110))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110110))
      begin
        rob__27_com_2 = soc2.core.rob.rob_uop__27_br_mask;
        rob__27_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__27_com_2 = 12'h0;
        rob__27_uncom_2 = soc2.core.rob.rob_uop__27_br_mask;
      end
    end
  end

  wire [11:0] rob__28_com_2;
  wire [11:0] rob__28_uncom_2;

  always @(*)
  begin
    rob__28_com_2 = 12'h0;
    rob__28_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b111000))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111000))
      begin
        rob__28_com_2 = soc2.core.rob.rob_uop__28_br_mask;
        rob__28_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__28_com_2 = 12'h0;
        rob__28_uncom_2 = soc2.core.rob.rob_uop__28_br_mask;
      end
    end
  end

  wire [11:0] rob__29_com_2;
  wire [11:0] rob__29_uncom_2;

  always @(*)
  begin
    rob__29_com_2 = 12'h0;
    rob__29_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b111010))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111010))
      begin
        rob__29_com_2 = soc2.core.rob.rob_uop__29_br_mask;
        rob__29_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__29_com_2 = 12'h0;
        rob__29_uncom_2 = soc2.core.rob.rob_uop__29_br_mask;
      end
    end
  end

  wire [11:0] rob__30_com_2;
  wire [11:0] rob__30_uncom_2;

  always @(*)
  begin
    rob__30_com_2 = 12'h0;
    rob__30_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b111100))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111100))
      begin
        rob__30_com_2 = soc2.core.rob.rob_uop__30_br_mask;
        rob__30_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__30_com_2 = 12'h0;
        rob__30_uncom_2 = soc2.core.rob.rob_uop__30_br_mask;
      end
    end
  end

  wire [11:0] rob__31_com_2;
  wire [11:0] rob__31_uncom_2;

  always @(*)
  begin
    rob__31_com_2 = 12'h0;
    rob__31_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b111110))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111110))
      begin
        rob__31_com_2 = soc2.core.rob.rob_uop__31_br_mask;
        rob__31_uncom_2 = 12'hfff;
      end
      else
      begin
        rob__31_com_2 = 12'h0;
        rob__31_uncom_2 = soc2.core.rob.rob_uop__31_br_mask;
      end
    end
  end

  wire [11:0] rob_1_0_com_2;
  wire [11:0] rob_1_0_uncom_2;

  always @(*)
  begin
    rob_1_0_com_2 = 12'h0;
    rob_1_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b000001))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000001))
      begin
        rob_1_0_com_2 = soc2.core.rob.rob_uop_1_0_br_mask;
        rob_1_0_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_0_com_2 = 12'h0;
        rob_1_0_uncom_2 = soc2.core.rob.rob_uop_1_0_br_mask;
      end
    end
  end

  wire [11:0] rob_1_1_com_2;
  wire [11:0] rob_1_1_uncom_2;

  always @(*)
  begin
    rob_1_1_com_2 = 12'h0;
    rob_1_1_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b000011))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000011))
      begin
        rob_1_1_com_2 = soc2.core.rob.rob_uop_1_1_br_mask;
        rob_1_1_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_1_com_2 = 12'h0;
        rob_1_1_uncom_2 = soc2.core.rob.rob_uop_1_1_br_mask;
      end
    end
  end

  wire [11:0] rob_1_2_com_2;
  wire [11:0] rob_1_2_uncom_2;

  always @(*)
  begin
    rob_1_2_com_2 = 12'h0;
    rob_1_2_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b000101))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000101))
      begin
        rob_1_2_com_2 = soc2.core.rob.rob_uop_1_2_br_mask;
        rob_1_2_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_2_com_2 = 12'h0;
        rob_1_2_uncom_2 = soc2.core.rob.rob_uop_1_2_br_mask;
      end
    end
  end

  wire [11:0] rob_1_3_com_2;
  wire [11:0] rob_1_3_uncom_2;

  always @(*)
  begin
    rob_1_3_com_2 = 12'h0;
    rob_1_3_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b000111))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b000111))
      begin
        rob_1_3_com_2 = soc2.core.rob.rob_uop_1_3_br_mask;
        rob_1_3_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_3_com_2 = 12'h0;
        rob_1_3_uncom_2 = soc2.core.rob.rob_uop_1_3_br_mask;
      end
    end
  end

  wire [11:0] rob_1_4_com_2;
  wire [11:0] rob_1_4_uncom_2;

  always @(*)
  begin
    rob_1_4_com_2 = 12'h0;
    rob_1_4_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b001001))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001001))
      begin
        rob_1_4_com_2 = soc2.core.rob.rob_uop_1_4_br_mask;
        rob_1_4_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_4_com_2 = 12'h0;
        rob_1_4_uncom_2 = soc2.core.rob.rob_uop_1_4_br_mask;
      end
    end
  end

  wire [11:0] rob_1_5_com_2;
  wire [11:0] rob_1_5_uncom_2;

  always @(*)
  begin
    rob_1_5_com_2 = 12'h0;
    rob_1_5_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b001011))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001011))
      begin
        rob_1_5_com_2 = soc2.core.rob.rob_uop_1_5_br_mask;
        rob_1_5_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_5_com_2 = 12'h0;
        rob_1_5_uncom_2 = soc2.core.rob.rob_uop_1_5_br_mask;
      end
    end
  end

  wire [11:0] rob_1_6_com_2;
  wire [11:0] rob_1_6_uncom_2;

  always @(*)
  begin
    rob_1_6_com_2 = 12'h0;
    rob_1_6_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b001101))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001101))
      begin
        rob_1_6_com_2 = soc2.core.rob.rob_uop_1_6_br_mask;
        rob_1_6_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_6_com_2 = 12'h0;
        rob_1_6_uncom_2 = soc2.core.rob.rob_uop_1_6_br_mask;
      end
    end
  end

  wire [11:0] rob_1_7_com_2;
  wire [11:0] rob_1_7_uncom_2;

  always @(*)
  begin
    rob_1_7_com_2 = 12'h0;
    rob_1_7_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b001111))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b001111))
      begin
        rob_1_7_com_2 = soc2.core.rob.rob_uop_1_7_br_mask;
        rob_1_7_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_7_com_2 = 12'h0;
        rob_1_7_uncom_2 = soc2.core.rob.rob_uop_1_7_br_mask;
      end
    end
  end

  wire [11:0] rob_1_8_com_2;
  wire [11:0] rob_1_8_uncom_2;

  always @(*)
  begin
    rob_1_8_com_2 = 12'h0;
    rob_1_8_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b010001))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010001))
      begin
        rob_1_8_com_2 = soc2.core.rob.rob_uop_1_8_br_mask;
        rob_1_8_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_8_com_2 = 12'h0;
        rob_1_8_uncom_2 = soc2.core.rob.rob_uop_1_8_br_mask;
      end
    end
  end

  wire [11:0] rob_1_9_com_2;
  wire [11:0] rob_1_9_uncom_2;

  always @(*)
  begin
    rob_1_9_com_2 = 12'h0;
    rob_1_9_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b010011))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010011))
      begin
        rob_1_9_com_2 = soc2.core.rob.rob_uop_1_9_br_mask;
        rob_1_9_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_9_com_2 = 12'h0;
        rob_1_9_uncom_2 = soc2.core.rob.rob_uop_1_9_br_mask;
      end
    end
  end

  wire [11:0] rob_1_10_com_2;
  wire [11:0] rob_1_10_uncom_2;

  always @(*)
  begin
    rob_1_10_com_2 = 12'h0;
    rob_1_10_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b010101))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010101))
      begin
        rob_1_10_com_2 = soc2.core.rob.rob_uop_1_10_br_mask;
        rob_1_10_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_10_com_2 = 12'h0;
        rob_1_10_uncom_2 = soc2.core.rob.rob_uop_1_10_br_mask;
      end
    end
  end

  wire [11:0] rob_1_11_com_2;
  wire [11:0] rob_1_11_uncom_2;

  always @(*)
  begin
    rob_1_11_com_2 = 12'h0;
    rob_1_11_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b010111))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b010111))
      begin
        rob_1_11_com_2 = soc2.core.rob.rob_uop_1_11_br_mask;
        rob_1_11_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_11_com_2 = 12'h0;
        rob_1_11_uncom_2 = soc2.core.rob.rob_uop_1_11_br_mask;
      end
    end
  end

  wire [11:0] rob_1_12_com_2;
  wire [11:0] rob_1_12_uncom_2;

  always @(*)
  begin
    rob_1_12_com_2 = 12'h0;
    rob_1_12_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b011001))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011001))
      begin
        rob_1_12_com_2 = soc2.core.rob.rob_uop_1_12_br_mask;
        rob_1_12_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_12_com_2 = 12'h0;
        rob_1_12_uncom_2 = soc2.core.rob.rob_uop_1_12_br_mask;
      end
    end
  end

  wire [11:0] rob_1_13_com_2;
  wire [11:0] rob_1_13_uncom_2;

  always @(*)
  begin
    rob_1_13_com_2 = 12'h0;
    rob_1_13_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b011011))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011011))
      begin
        rob_1_13_com_2 = soc2.core.rob.rob_uop_1_13_br_mask;
        rob_1_13_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_13_com_2 = 12'h0;
        rob_1_13_uncom_2 = soc2.core.rob.rob_uop_1_13_br_mask;
      end
    end
  end

  wire [11:0] rob_1_14_com_2;
  wire [11:0] rob_1_14_uncom_2;

  always @(*)
  begin
    rob_1_14_com_2 = 12'h0;
    rob_1_14_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b011101))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011101))
      begin
        rob_1_14_com_2 = soc2.core.rob.rob_uop_1_14_br_mask;
        rob_1_14_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_14_com_2 = 12'h0;
        rob_1_14_uncom_2 = soc2.core.rob.rob_uop_1_14_br_mask;
      end
    end
  end

  wire [11:0] rob_1_15_com_2;
  wire [11:0] rob_1_15_uncom_2;

  always @(*)
  begin
    rob_1_15_com_2 = 12'h0;
    rob_1_15_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b011111))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b011111))
      begin
        rob_1_15_com_2 = soc2.core.rob.rob_uop_1_15_br_mask;
        rob_1_15_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_15_com_2 = 12'h0;
        rob_1_15_uncom_2 = soc2.core.rob.rob_uop_1_15_br_mask;
      end
    end
  end

  wire [11:0] rob_1_16_com_2;
  wire [11:0] rob_1_16_uncom_2;

  always @(*)
  begin
    rob_1_16_com_2 = 12'h0;
    rob_1_16_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b100001))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100001))
      begin
        rob_1_16_com_2 = soc2.core.rob.rob_uop_1_16_br_mask;
        rob_1_16_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_16_com_2 = 12'h0;
        rob_1_16_uncom_2 = soc2.core.rob.rob_uop_1_16_br_mask;
      end
    end
  end

  wire [11:0] rob_1_17_com_2;
  wire [11:0] rob_1_17_uncom_2;

  always @(*)
  begin
    rob_1_17_com_2 = 12'h0;
    rob_1_17_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b100011))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100011))
      begin
        rob_1_17_com_2 = soc2.core.rob.rob_uop_1_17_br_mask;
        rob_1_17_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_17_com_2 = 12'h0;
        rob_1_17_uncom_2 = soc2.core.rob.rob_uop_1_17_br_mask;
      end
    end
  end

  wire [11:0] rob_1_18_com_2;
  wire [11:0] rob_1_18_uncom_2;

  always @(*)
  begin
    rob_1_18_com_2 = 12'h0;
    rob_1_18_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b100101))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100101))
      begin
        rob_1_18_com_2 = soc2.core.rob.rob_uop_1_18_br_mask;
        rob_1_18_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_18_com_2 = 12'h0;
        rob_1_18_uncom_2 = soc2.core.rob.rob_uop_1_18_br_mask;
      end
    end
  end

  wire [11:0] rob_1_19_com_2;
  wire [11:0] rob_1_19_uncom_2;

  always @(*)
  begin
    rob_1_19_com_2 = 12'h0;
    rob_1_19_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b100111))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b100111))
      begin
        rob_1_19_com_2 = soc2.core.rob.rob_uop_1_19_br_mask;
        rob_1_19_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_19_com_2 = 12'h0;
        rob_1_19_uncom_2 = soc2.core.rob.rob_uop_1_19_br_mask;
      end
    end
  end

  wire [11:0] rob_1_20_com_2;
  wire [11:0] rob_1_20_uncom_2;

  always @(*)
  begin
    rob_1_20_com_2 = 12'h0;
    rob_1_20_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b101001))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101001))
      begin
        rob_1_20_com_2 = soc2.core.rob.rob_uop_1_20_br_mask;
        rob_1_20_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_20_com_2 = 12'h0;
        rob_1_20_uncom_2 = soc2.core.rob.rob_uop_1_20_br_mask;
      end
    end
  end

  wire [11:0] rob_1_21_com_2;
  wire [11:0] rob_1_21_uncom_2;

  always @(*)
  begin
    rob_1_21_com_2 = 12'h0;
    rob_1_21_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b101011))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101011))
      begin
        rob_1_21_com_2 = soc2.core.rob.rob_uop_1_21_br_mask;
        rob_1_21_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_21_com_2 = 12'h0;
        rob_1_21_uncom_2 = soc2.core.rob.rob_uop_1_21_br_mask;
      end
    end
  end

  wire [11:0] rob_1_22_com_2;
  wire [11:0] rob_1_22_uncom_2;

  always @(*)
  begin
    rob_1_22_com_2 = 12'h0;
    rob_1_22_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b101101))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101101))
      begin
        rob_1_22_com_2 = soc2.core.rob.rob_uop_1_22_br_mask;
        rob_1_22_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_22_com_2 = 12'h0;
        rob_1_22_uncom_2 = soc2.core.rob.rob_uop_1_22_br_mask;
      end
    end
  end

  wire [11:0] rob_1_23_com_2;
  wire [11:0] rob_1_23_uncom_2;

  always @(*)
  begin
    rob_1_23_com_2 = 12'h0;
    rob_1_23_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b101111))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b101111))
      begin
        rob_1_23_com_2 = soc2.core.rob.rob_uop_1_23_br_mask;
        rob_1_23_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_23_com_2 = 12'h0;
        rob_1_23_uncom_2 = soc2.core.rob.rob_uop_1_23_br_mask;
      end
    end
  end

  wire [11:0] rob_1_24_com_2;
  wire [11:0] rob_1_24_uncom_2;

  always @(*)
  begin
    rob_1_24_com_2 = 12'h0;
    rob_1_24_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b110001))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110001))
      begin
        rob_1_24_com_2 = soc2.core.rob.rob_uop_1_24_br_mask;
        rob_1_24_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_24_com_2 = 12'h0;
        rob_1_24_uncom_2 = soc2.core.rob.rob_uop_1_24_br_mask;
      end
    end
  end

  wire [11:0] rob_1_25_com_2;
  wire [11:0] rob_1_25_uncom_2;

  always @(*)
  begin
    rob_1_25_com_2 = 12'h0;
    rob_1_25_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b110011))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110011))
      begin
        rob_1_25_com_2 = soc2.core.rob.rob_uop_1_25_br_mask;
        rob_1_25_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_25_com_2 = 12'h0;
        rob_1_25_uncom_2 = soc2.core.rob.rob_uop_1_25_br_mask;
      end
    end
  end

  wire [11:0] rob_1_26_com_2;
  wire [11:0] rob_1_26_uncom_2;

  always @(*)
  begin
    rob_1_26_com_2 = 12'h0;
    rob_1_26_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b110101))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110101))
      begin
        rob_1_26_com_2 = soc2.core.rob.rob_uop_1_26_br_mask;
        rob_1_26_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_26_com_2 = 12'h0;
        rob_1_26_uncom_2 = soc2.core.rob.rob_uop_1_26_br_mask;
      end
    end
  end

  wire [11:0] rob_1_27_com_2;
  wire [11:0] rob_1_27_uncom_2;

  always @(*)
  begin
    rob_1_27_com_2 = 12'h0;
    rob_1_27_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b110111))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b110111))
      begin
        rob_1_27_com_2 = soc2.core.rob.rob_uop_1_27_br_mask;
        rob_1_27_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_27_com_2 = 12'h0;
        rob_1_27_uncom_2 = soc2.core.rob.rob_uop_1_27_br_mask;
      end
    end
  end

  wire [11:0] rob_1_28_com_2;
  wire [11:0] rob_1_28_uncom_2;

  always @(*)
  begin
    rob_1_28_com_2 = 12'h0;
    rob_1_28_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b111001))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111001))
      begin
        rob_1_28_com_2 = soc2.core.rob.rob_uop_1_28_br_mask;
        rob_1_28_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_28_com_2 = 12'h0;
        rob_1_28_uncom_2 = soc2.core.rob.rob_uop_1_28_br_mask;
      end
    end
  end

  wire [11:0] rob_1_29_com_2;
  wire [11:0] rob_1_29_uncom_2;

  always @(*)
  begin
    rob_1_29_com_2 = 12'h0;
    rob_1_29_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b111011))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111011))
      begin
        rob_1_29_com_2 = soc2.core.rob.rob_uop_1_29_br_mask;
        rob_1_29_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_29_com_2 = 12'h0;
        rob_1_29_uncom_2 = soc2.core.rob.rob_uop_1_29_br_mask;
      end
    end
  end

  wire [11:0] rob_1_30_com_2;
  wire [11:0] rob_1_30_uncom_2;

  always @(*)
  begin
    rob_1_30_com_2 = 12'h0;
    rob_1_30_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b111101))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111101))
      begin
        rob_1_30_com_2 = soc2.core.rob.rob_uop_1_30_br_mask;
        rob_1_30_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_30_com_2 = 12'h0;
        rob_1_30_uncom_2 = soc2.core.rob.rob_uop_1_30_br_mask;
      end
    end
  end

  wire [11:0] rob_1_31_com_2;
  wire [11:0] rob_1_31_uncom_2;

  always @(*)
  begin
    rob_1_31_com_2 = 12'h0;
    rob_1_31_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(6'b111111))
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, 6'b111111))
      begin
        rob_1_31_com_2 = soc2.core.rob.rob_uop_1_31_br_mask;
        rob_1_31_uncom_2 = 12'hfff;
      end
      else
      begin
        rob_1_31_com_2 = 12'h0;
        rob_1_31_uncom_2 = soc2.core.rob.rob_uop_1_31_br_mask;
      end
    end
  end

  wire [11:0] lsu_clr_bsy_brmask_0_com_2;
  wire [11:0] lsu_clr_bsy_brmask_0_uncom_2;

  always @(*)
  begin
    lsu_clr_bsy_brmask_0_com_2 = 12'h0;
    lsu_clr_bsy_brmask_0_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.clr_bsy_rob_idx_0) && soc2.lsu.clr_bsy_valid_0)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.clr_bsy_rob_idx_0))
      begin
        lsu_clr_bsy_brmask_0_com_2 = soc2.lsu.clr_bsy_brmask_0;
        lsu_clr_bsy_brmask_0_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_clr_bsy_brmask_0_com_2 = 12'h0;
        lsu_clr_bsy_brmask_0_uncom_2 = soc2.lsu.clr_bsy_brmask_0;
      end
    end
  end

  wire [11:0] lsu_r_xcpt_com_2;
  wire [11:0] lsu_r_xcpt_uncom_2;

  always @(*)
  begin
    lsu_r_xcpt_com_2 = 12'h0;
    lsu_r_xcpt_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(soc2.lsu.r_xcpt_uop_rob_idx) && soc2.lsu.r_xcpt_valid)
    begin
      if (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.r_xcpt_uop_rob_idx))
      begin
        lsu_r_xcpt_com_2 = soc2.lsu.r_xcpt_uop_br_mask;
        lsu_r_xcpt_uncom_2 = 12'hfff;
      end
      else
      begin
        lsu_r_xcpt_com_2 = 12'h0;
        lsu_r_xcpt_uncom_2 = soc2.lsu.r_xcpt_uop_br_mask;
      end
    end
  end

  //bookkeeping buffers without explicit rob_idx
  //check if loadqueue/storequeue are used and get ROB ID from ldq_idx/stq_idx

  wire [11:0] respq_uops_0_ldq_com_2;
  wire [11:0] respq_uops_0_ldq_uncom_2;

  always @(*)
  begin
    respq_uops_0_ldq_com_2 = 12'h0;
    respq_uops_0_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_0_ldq_idx]) && soc2.dcache.mshrs.respq.valids_0)
    begin
      if(soc2.dcache.mshrs.respq.uops_0_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_0_ldq_idx]))
        begin
          respq_uops_0_ldq_com_2 = soc2.dcache.mshrs.respq.uops_0_br_mask;
          respq_uops_0_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          respq_uops_0_ldq_com_2 = 12'h0;
          respq_uops_0_ldq_uncom_2 = soc2.dcache.mshrs.respq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_1_ldq_com_2;
  wire [11:0] respq_uops_1_ldq_uncom_2;

  always @(*)
  begin
    respq_uops_1_ldq_com_2 = 12'h0;
    respq_uops_1_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_1_ldq_idx]) && soc2.dcache.mshrs.respq.valids_1)
    begin
      if(soc2.dcache.mshrs.respq.uops_1_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_1_ldq_idx]))
        begin
          respq_uops_1_ldq_com_2 = soc2.dcache.mshrs.respq.uops_1_br_mask;
          respq_uops_1_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          respq_uops_1_ldq_com_2 = 12'h0;
          respq_uops_1_ldq_uncom_2 = soc2.dcache.mshrs.respq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_2_ldq_com_2;
  wire [11:0] respq_uops_2_ldq_uncom_2;

  always @(*)
  begin
    respq_uops_2_ldq_com_2 = 12'h0;
    respq_uops_2_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_2_ldq_idx]) && soc2.dcache.mshrs.respq.valids_2)
    begin
      if(soc2.dcache.mshrs.respq.uops_2_uses_ldq == 1'b1)
      begin
      if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_2_ldq_idx]))
        begin
          respq_uops_2_ldq_com_2 = soc2.dcache.mshrs.respq.uops_2_br_mask;
          respq_uops_2_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          respq_uops_2_ldq_com_2 = 12'h0;
          respq_uops_2_ldq_uncom_2 = soc2.dcache.mshrs.respq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_3_ldq_com_2;
  wire [11:0] respq_uops_3_ldq_uncom_2;

  always @(*)
  begin
    respq_uops_3_ldq_com_2 = 12'h0;
    respq_uops_3_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_3_ldq_idx]) && soc2.dcache.mshrs.respq.valids_3)
    begin
      if(soc2.dcache.mshrs.respq.uops_3_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_3_ldq_idx]))
        begin
          respq_uops_3_ldq_com_2 = soc2.dcache.mshrs.respq.uops_3_br_mask;
          respq_uops_3_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          respq_uops_3_ldq_com_2 = 12'h0;
          respq_uops_3_ldq_uncom_2 = soc2.dcache.mshrs.respq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_0_stq_com_2;
  wire [11:0] respq_uops_0_stq_uncom_2;

  always @(*)
  begin
    respq_uops_0_stq_com_2 = 12'h0;
    respq_uops_0_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_0_stq_idx]) && soc2.dcache.mshrs.respq.valids_0 && !(soc2.dcache.mshrs.respq.uops_0_uses_stq && stq_committed_2[soc2.dcache.mshrs.respq.uops_0_stq_idx]))
    begin
      if(soc2.dcache.mshrs.respq.uops_0_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_0_stq_idx]))
        begin
          respq_uops_0_stq_com_2 = soc2.dcache.mshrs.respq.uops_0_br_mask;
          respq_uops_0_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          respq_uops_0_stq_com_2 = 12'h0;
          respq_uops_0_stq_uncom_2 = soc2.dcache.mshrs.respq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_1_stq_com_2;
  wire [11:0] respq_uops_1_stq_uncom_2;

  always @(*)
  begin
    respq_uops_1_stq_com_2 = 12'h0;
    respq_uops_1_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_1_stq_idx]) && soc2.dcache.mshrs.respq.valids_1 && !(soc2.dcache.mshrs.respq.uops_1_uses_stq && stq_committed_2[soc2.dcache.mshrs.respq.uops_1_stq_idx]))
    begin
      if(soc2.dcache.mshrs.respq.uops_1_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_1_stq_idx]))
        begin
          respq_uops_1_stq_com_2 = soc2.dcache.mshrs.respq.uops_1_br_mask;
          respq_uops_1_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          respq_uops_1_stq_com_2 = 12'h0;
          respq_uops_1_stq_uncom_2 = soc2.dcache.mshrs.respq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_2_stq_com_2;
  wire [11:0] respq_uops_2_stq_uncom_2;

  always @(*)
  begin
    respq_uops_2_stq_com_2 = 12'h0;
    respq_uops_2_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_2_stq_idx]) && soc2.dcache.mshrs.respq.valids_2 && !(soc2.dcache.mshrs.respq.uops_2_uses_stq && stq_committed_2[soc2.dcache.mshrs.respq.uops_2_stq_idx]))
    begin
      if(soc2.dcache.mshrs.respq.uops_2_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_2_stq_idx]))
        begin
          respq_uops_2_stq_com_2 = soc2.dcache.mshrs.respq.uops_2_br_mask;
          respq_uops_2_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          respq_uops_2_stq_com_2 = 12'h0;
          respq_uops_2_stq_uncom_2 = soc2.dcache.mshrs.respq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] respq_uops_3_stq_com_2;
  wire [11:0] respq_uops_3_stq_uncom_2;

  always @(*)
  begin
    respq_uops_3_stq_com_2 = 12'h0;
    respq_uops_3_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_3_stq_idx]) && soc2.dcache.mshrs.respq.valids_3 && !(soc2.dcache.mshrs.respq.uops_3_uses_stq && stq_committed_2[soc2.dcache.mshrs.respq.uops_3_stq_idx]))
    begin
      if(soc2.dcache.mshrs.respq.uops_3_uses_stq == 1'b1)
      begin
      if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_3_stq_idx]))
        begin
          respq_uops_3_stq_com_2 = soc2.dcache.mshrs.respq.uops_3_br_mask;
          respq_uops_3_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          respq_uops_3_stq_com_2 = 12'h0;
          respq_uops_3_stq_uncom_2 = soc2.dcache.mshrs.respq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mmios_0_ldq_com_2;
  wire [11:0] mmios_0_ldq_uncom_2;

  always @(*)
  begin
    mmios_0_ldq_com_2 = 12'h0;
    mmios_0_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mmios_0.req_uop_ldq_idx]) && soc2.dcache.mshrs.mmios_0.state != 2'b0)
    begin
      if(soc2.dcache.mshrs.mmios_0.req_uop_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mmios_0.req_uop_ldq_idx]))
        begin
          mmios_0_ldq_com_2 = soc2.dcache.mshrs.mmios_0.req_uop_br_mask;
          mmios_0_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mmios_0_ldq_com_2 = 12'h0;
          mmios_0_ldq_uncom_2 = soc2.dcache.mshrs.mmios_0.req_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] mmios_0_stq_com_2;
  wire [11:0] mmios_0_stq_uncom_2;

  always @(*)
  begin
    mmios_0_stq_com_2 = 12'h0;
    mmios_0_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mmios_0.req_uop_stq_idx]) && soc2.dcache.mshrs.mmios_0.state != 2'b0)
    begin
      if((soc2.dcache.mshrs.mmios_0.req_uop_uses_stq == 1'b1) && !stq_committed_2[soc2.dcache.mshrs.mmios_0.req_uop_stq_idx])
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mmios_0.req_uop_stq_idx]))
        begin
          mmios_0_stq_com_2 = soc2.dcache.mshrs.mmios_0.req_uop_br_mask;
          mmios_0_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mmios_0_stq_com_2 = 12'h0;
          mmios_0_stq_uncom_2 = soc2.dcache.mshrs.mmios_0.req_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_0_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_0_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_0_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_0_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_0_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_0)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_0_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_0_ldq_idx]))
        begin
          mshrs_0_rpq_uops_0_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask;
          mshrs_0_rpq_uops_0_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_0_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_0_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_1_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_1_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_1_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_1_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_1_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_1)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_1_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_1_ldq_idx]))
        begin
          mshrs_0_rpq_uops_1_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask;
          mshrs_0_rpq_uops_1_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_1_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_1_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_2_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_2_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_2_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_2_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_2_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_2)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_2_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_2_ldq_idx]))
        begin
          mshrs_0_rpq_uops_2_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask;
          mshrs_0_rpq_uops_2_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_2_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_2_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_3_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_3_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_3_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_3_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_3_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_3)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_3_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_3_ldq_idx]))
        begin
          mshrs_0_rpq_uops_3_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask;
          mshrs_0_rpq_uops_3_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_3_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_3_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_4_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_4_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_4_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_4_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_4_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_4)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_4_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_4_ldq_idx]))
        begin
          mshrs_0_rpq_uops_4_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask;
          mshrs_0_rpq_uops_4_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_4_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_4_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_5_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_5_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_5_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_5_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_5_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_5)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_5_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_5_ldq_idx]))
        begin
          mshrs_0_rpq_uops_5_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask;
          mshrs_0_rpq_uops_5_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_5_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_5_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_6_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_6_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_6_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_6_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_6_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_6)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_6_uses_ldq == 1'b1)
      begin
      if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_6_ldq_idx]))
        begin
          mshrs_0_rpq_uops_6_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask;
          mshrs_0_rpq_uops_6_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_6_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_6_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_7_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_7_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_7_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_7_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_7_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_7)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_7_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_7_ldq_idx]))
        begin
          mshrs_0_rpq_uops_7_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask;
          mshrs_0_rpq_uops_7_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_7_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_7_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_8_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_8_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_8_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_8_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_8_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_8)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_8_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_8_ldq_idx]))
        begin
          mshrs_0_rpq_uops_8_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask;
          mshrs_0_rpq_uops_8_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_8_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_8_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_9_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_9_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_9_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_9_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_9_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_9)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_9_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_9_ldq_idx]))
        begin
          mshrs_0_rpq_uops_9_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask;
          mshrs_0_rpq_uops_9_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_9_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_9_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_10_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_10_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_10_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_10_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_10_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_10)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_10_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_10_ldq_idx]))
        begin
          mshrs_0_rpq_uops_10_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask;
          mshrs_0_rpq_uops_10_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_10_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_10_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_11_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_11_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_11_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_11_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_11_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_11)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_11_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_11_ldq_idx]))
        begin
          mshrs_0_rpq_uops_11_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask;
          mshrs_0_rpq_uops_11_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_11_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_11_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_12_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_12_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_12_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_12_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_12_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_12)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_12_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_12_ldq_idx]))
        begin
          mshrs_0_rpq_uops_12_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask;
          mshrs_0_rpq_uops_12_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_12_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_12_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_13_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_13_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_13_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_13_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_13_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_13)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_13_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_13_ldq_idx]))
        begin
          mshrs_0_rpq_uops_13_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask;
          mshrs_0_rpq_uops_13_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_13_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_13_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_14_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_14_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_14_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_14_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_14_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_14)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_14_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_14_ldq_idx]))
        begin
          mshrs_0_rpq_uops_14_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask;
          mshrs_0_rpq_uops_14_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_14_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_14_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_15_ldq_com_2;
  wire [11:0] mshrs_0_rpq_uops_15_ldq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_15_ldq_com_2 = 12'h0;
    mshrs_0_rpq_uops_15_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_15_ldq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_15)
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_15_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_15_ldq_idx]))
        begin
          mshrs_0_rpq_uops_15_ldq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask;
          mshrs_0_rpq_uops_15_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_15_ldq_com_2 = 12'h0;
          mshrs_0_rpq_uops_15_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask;
        end
      end
    end
  end


  wire [11:0] mshrs_0_rpq_uops_0_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_0_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_0_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_0_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_0 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_0_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx]))
        begin
          mshrs_0_rpq_uops_0_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask;
          mshrs_0_rpq_uops_0_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_0_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_0_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_1_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_1_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_1_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_1_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_1 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_1_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx]))
        begin
          mshrs_0_rpq_uops_1_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask;
          mshrs_0_rpq_uops_1_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_1_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_1_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_2_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_2_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_2_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_2_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_2 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_2_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx]))
        begin
          mshrs_0_rpq_uops_2_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask;
          mshrs_0_rpq_uops_2_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_2_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_2_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_3_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_3_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_3_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_3_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_3 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_3_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx]))
        begin
          mshrs_0_rpq_uops_3_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask;
          mshrs_0_rpq_uops_3_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_3_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_3_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_4_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_4_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_4_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_4_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_4 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_4_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx]))
        begin
          mshrs_0_rpq_uops_4_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask;
          mshrs_0_rpq_uops_4_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_4_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_4_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_5_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_5_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_5_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_5_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_5 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_5_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx]))
        begin
          mshrs_0_rpq_uops_5_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask;
          mshrs_0_rpq_uops_5_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_5_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_5_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_6_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_6_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_6_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_6_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_6 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_6_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx]))
        begin
          mshrs_0_rpq_uops_6_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask;
          mshrs_0_rpq_uops_6_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_6_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_6_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_7_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_7_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_7_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_7_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_7 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_7_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx]))
        begin
          mshrs_0_rpq_uops_7_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask;
          mshrs_0_rpq_uops_7_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_7_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_7_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_8_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_8_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_8_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_8_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_8 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_8_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx]))
        begin
          mshrs_0_rpq_uops_8_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask;
          mshrs_0_rpq_uops_8_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_8_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_8_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_9_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_9_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_9_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_9_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_9 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_9_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx]))
        begin
          mshrs_0_rpq_uops_9_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask;
          mshrs_0_rpq_uops_9_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_9_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_9_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_10_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_10_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_10_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_10_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_10 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_10_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx]))
        begin
          mshrs_0_rpq_uops_10_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask;
          mshrs_0_rpq_uops_10_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_10_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_10_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_11_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_11_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_11_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_11_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_11 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_11_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx]))
        begin
          mshrs_0_rpq_uops_11_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask;
          mshrs_0_rpq_uops_11_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_11_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_11_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_12_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_12_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_12_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_12_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_12 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_12_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx]))
        begin
          mshrs_0_rpq_uops_12_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask;
          mshrs_0_rpq_uops_12_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_12_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_12_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_13_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_13_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_13_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_13_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_13 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_13_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx]))
        begin
          mshrs_0_rpq_uops_13_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask;
          mshrs_0_rpq_uops_13_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_13_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_13_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_14_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_14_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_14_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_14_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_14 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_14_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx]))
        begin
          mshrs_0_rpq_uops_14_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask;
          mshrs_0_rpq_uops_14_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_14_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_14_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_0_rpq_uops_15_stq_com_2;
  wire [11:0] mshrs_0_rpq_uops_15_stq_uncom_2;

  always @(*)
  begin
    mshrs_0_rpq_uops_15_stq_com_2 = 12'h0;
    mshrs_0_rpq_uops_15_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx]) && soc2.dcache.mshrs.mshrs_0.rpq.valids_15 && !stq_committed_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_0.rpq.uops_15_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx]))
        begin
          mshrs_0_rpq_uops_15_stq_com_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask;
          mshrs_0_rpq_uops_15_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_0_rpq_uops_15_stq_com_2 = 12'h0;
          mshrs_0_rpq_uops_15_stq_uncom_2 = soc2.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_0_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_0_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_0_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_0_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_0_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_0)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_0_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_0_ldq_idx]))
        begin
          mshrs_1_rpq_uops_0_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask;
          mshrs_1_rpq_uops_0_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_0_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_0_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_1_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_1_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_1_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_1_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_1_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_1)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_1_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_1_ldq_idx]))
        begin
          mshrs_1_rpq_uops_1_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask;
          mshrs_1_rpq_uops_1_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_0_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_0_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_2_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_2_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_2_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_2_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_2_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_2)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_2_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_2_ldq_idx]))
        begin
          mshrs_1_rpq_uops_2_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask;
          mshrs_1_rpq_uops_2_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_2_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_2_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_3_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_3_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_3_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_3_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_3_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_3)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_3_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_3_ldq_idx]))
        begin
          mshrs_1_rpq_uops_3_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask;
          mshrs_1_rpq_uops_3_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_3_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_3_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_4_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_4_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_4_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_4_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_4_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_4)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_4_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_4_ldq_idx]))
        begin
          mshrs_1_rpq_uops_4_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask;
          mshrs_1_rpq_uops_4_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_4_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_4_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_5_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_5_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_5_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_5_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_5_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_5)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_5_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_5_ldq_idx]))
        begin
          mshrs_1_rpq_uops_5_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask;
          mshrs_1_rpq_uops_5_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_5_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_5_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_6_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_6_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_6_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_6_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_6_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_6)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_6_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_6_ldq_idx]))
        begin
          mshrs_1_rpq_uops_6_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask;
          mshrs_1_rpq_uops_6_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_6_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_6_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_7_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_7_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_7_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_7_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_7_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_7)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_7_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_7_ldq_idx]))
        begin
          mshrs_1_rpq_uops_7_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask;
          mshrs_1_rpq_uops_7_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_7_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_7_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_8_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_8_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_8_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_8_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_8_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_8)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_8_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_8_ldq_idx]))
        begin
          mshrs_1_rpq_uops_8_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask;
          mshrs_1_rpq_uops_8_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_8_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_8_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_9_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_9_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_9_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_9_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_9_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_9)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_9_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_9_ldq_idx]))
        begin
          mshrs_1_rpq_uops_9_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask;
          mshrs_1_rpq_uops_9_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_9_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_9_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_10_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_10_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_10_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_10_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_10_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_10)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_10_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_10_ldq_idx]))
        begin
          mshrs_1_rpq_uops_10_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask;
          mshrs_1_rpq_uops_10_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_10_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_10_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_11_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_11_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_11_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_11_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_11_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_11)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_11_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_11_ldq_idx]))
        begin
          mshrs_1_rpq_uops_11_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask;
          mshrs_1_rpq_uops_11_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_11_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_11_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_12_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_12_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_12_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_12_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_12_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_12)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_12_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_12_ldq_idx]))
        begin
          mshrs_1_rpq_uops_12_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask;
          mshrs_1_rpq_uops_12_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_12_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_12_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_13_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_13_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_13_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_13_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_13_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_13)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_13_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_13_ldq_idx]))
        begin
          mshrs_1_rpq_uops_13_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask;
          mshrs_1_rpq_uops_13_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_13_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_13_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_14_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_14_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_14_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_14_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_14_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_14)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_14_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_14_ldq_idx]))
        begin
          mshrs_1_rpq_uops_14_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask;
          mshrs_1_rpq_uops_14_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_14_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_14_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_15_ldq_com_2;
  wire [11:0] mshrs_1_rpq_uops_15_ldq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_15_ldq_com_2 = 12'h0;
    mshrs_1_rpq_uops_15_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_15_ldq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_15)
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_15_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_15_ldq_idx]))
        begin
          mshrs_1_rpq_uops_15_ldq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask;
          mshrs_1_rpq_uops_15_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_15_ldq_com_2 = 12'h0;
          mshrs_1_rpq_uops_15_ldq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask;
        end
      end
    end
  end


  wire [11:0] mshrs_1_rpq_uops_0_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_0_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_0_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_0_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_0 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_0_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx]))
        begin
          mshrs_1_rpq_uops_0_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask;
          mshrs_1_rpq_uops_0_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_0_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_0_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_1_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_1_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_1_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_1_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_1 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_1_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx]))
        begin
          mshrs_1_rpq_uops_1_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask;
          mshrs_1_rpq_uops_1_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_0_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_0_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_2_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_2_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_2_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_2_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_2 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_2_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx]))
        begin
          mshrs_1_rpq_uops_2_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask;
          mshrs_1_rpq_uops_2_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_2_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_2_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_3_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_3_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_3_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_3_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_3 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_3_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx]))
        begin
          mshrs_1_rpq_uops_3_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask;
          mshrs_1_rpq_uops_3_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_3_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_3_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_4_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_4_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_4_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_4_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_4 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_4_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx]))
        begin
          mshrs_1_rpq_uops_4_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask;
          mshrs_1_rpq_uops_4_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_4_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_4_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_5_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_5_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_5_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_5_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_5 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_5_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx]))
        begin
          mshrs_1_rpq_uops_5_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask;
          mshrs_1_rpq_uops_5_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_5_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_5_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_6_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_6_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_6_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_6_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_6 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_6_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx]))
        begin
          mshrs_1_rpq_uops_6_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask;
          mshrs_1_rpq_uops_6_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_6_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_6_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_7_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_7_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_7_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_7_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_7 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_7_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx]))
        begin
          mshrs_1_rpq_uops_7_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask;
          mshrs_1_rpq_uops_7_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_7_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_7_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_8_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_8_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_8_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_8_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_8 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_8_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx]))
        begin
          mshrs_1_rpq_uops_8_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask;
          mshrs_1_rpq_uops_8_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_8_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_8_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_9_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_9_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_9_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_9_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_9 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_9_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx]))
        begin
          mshrs_1_rpq_uops_9_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask;
          mshrs_1_rpq_uops_9_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_9_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_9_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_10_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_10_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_10_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_10_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_10 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_10_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx]))
        begin
          mshrs_1_rpq_uops_10_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask;
          mshrs_1_rpq_uops_10_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_10_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_10_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_11_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_11_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_11_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_11_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_11 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_11_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx]))
        begin
          mshrs_1_rpq_uops_11_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask;
          mshrs_1_rpq_uops_11_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_11_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_11_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_12_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_12_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_12_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_12_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_12 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_12_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx]))
        begin
          mshrs_1_rpq_uops_12_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask;
          mshrs_1_rpq_uops_12_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_12_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_12_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_13_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_13_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_13_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_13_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_13 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_13_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx]))
        begin
          mshrs_1_rpq_uops_13_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask;
          mshrs_1_rpq_uops_13_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_13_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_13_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_14_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_14_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_14_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_14_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_14 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_14_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx]))
        begin
          mshrs_1_rpq_uops_14_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask;
          mshrs_1_rpq_uops_14_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_14_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_14_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask;
        end
      end
    end
  end

  wire [11:0] mshrs_1_rpq_uops_15_stq_com_2;
  wire [11:0] mshrs_1_rpq_uops_15_stq_uncom_2;

  always @(*)
  begin
    mshrs_1_rpq_uops_15_stq_com_2 = 12'h0;
    mshrs_1_rpq_uops_15_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx]) && soc2.dcache.mshrs.mshrs_1.rpq.valids_15 && !stq_committed_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx])
    begin
      if(soc2.dcache.mshrs.mshrs_1.rpq.uops_15_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx]))
        begin
          mshrs_1_rpq_uops_15_stq_com_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask;
          mshrs_1_rpq_uops_15_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          mshrs_1_rpq_uops_15_stq_com_2 = 12'h0;
          mshrs_1_rpq_uops_15_stq_uncom_2 = soc2.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask;
        end
      end
    end
  end

  wire [11:0] dcache_s1_req_ldq_com_2;
  wire [11:0] dcache_s1_req_ldq_uncom_2;

  always @(*)
  begin
    dcache_s1_req_ldq_com_2 = 12'h0;
    dcache_s1_req_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.s1_req_0_uop_ldq_idx]) /*&& soc2.dcache.s1_valid_0*/)
    begin
      if(soc2.dcache.s1_req_0_uop_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.s1_req_0_uop_ldq_idx]))
        begin
          dcache_s1_req_ldq_com_2 = soc2.dcache.s1_req_0_uop_br_mask;
          dcache_s1_req_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          dcache_s1_req_ldq_com_2 = 12'h0;
          dcache_s1_req_ldq_uncom_2 = soc2.dcache.s1_req_0_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] dcache_s1_req_stq_com_2;
  wire [11:0] dcache_s1_req_stq_uncom_2;

  always @(*)
  begin
    dcache_s1_req_stq_com_2 = 12'h0;
    dcache_s1_req_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.s1_req_0_uop_stq_idx]) && /*soc2.dcache.s1_valid_0 &&*/ !stq_committed_2[soc2.dcache.s1_req_0_uop_stq_idx])
    begin
      if(soc2.dcache.s1_req_0_uop_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.s1_req_0_uop_stq_idx]))
        begin
          dcache_s1_req_stq_com_2 = soc2.dcache.s1_req_0_uop_br_mask;
          dcache_s1_req_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          dcache_s1_req_stq_com_2 = 12'h0;
          dcache_s1_req_stq_uncom_2 = soc2.dcache.s1_req_0_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] dcache_s2_req_ldq_com_2;
  wire [11:0] dcache_s2_req_ldq_uncom_2;

  always @(*)
  begin
    dcache_s2_req_ldq_com_2 = 12'h0;
    dcache_s2_req_ldq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(ldq_rob_idx_2[soc2.dcache.s2_req_0_uop_ldq_idx]) /*&& soc2.dcache.s2_valid_0*/)
    begin
      if(soc2.dcache.s2_req_0_uop_uses_ldq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.dcache.s2_req_0_uop_ldq_idx]))
        begin
          dcache_s2_req_ldq_com_2 = soc2.dcache.s2_req_0_uop_br_mask;
          dcache_s2_req_ldq_uncom_2 = 12'hfff;
        end
        else
        begin
          dcache_s2_req_ldq_com_2 = 12'h0;
          dcache_s2_req_ldq_uncom_2 = soc2.dcache.s2_req_0_uop_br_mask;
        end
      end
    end
  end

  wire [11:0] dcache_s2_req_stq_com_2;
  wire [11:0] dcache_s2_req_stq_uncom_2;

  always @(*)
  begin
    dcache_s2_req_stq_com_2 = 12'h0;
    dcache_s2_req_stq_uncom_2 = 12'hfff;
    if(isInBoundsROB_2(stq_rob_idx_2[soc2.dcache.s2_req_0_uop_stq_idx]) && /*soc2.dcache.s2_valid_0 && */!stq_committed_2[soc2.dcache.s2_req_0_uop_stq_idx])
    begin
      if(soc2.dcache.s2_req_0_uop_uses_stq == 1'b1)
      begin
        if(isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.dcache.s2_req_0_uop_stq_idx]))
        begin
          dcache_s2_req_stq_com_2 = soc2.dcache.s2_req_0_uop_br_mask;
          dcache_s2_req_stq_uncom_2 = 12'hfff;
        end
        else
        begin
          dcache_s2_req_stq_com_2 = 12'h0;
          dcache_s2_req_stq_uncom_2 = soc2.dcache.s2_req_0_uop_br_mask;
        end
      end
    end
  end

//*******************************************//
	wire [11:0] commitable_masks_2;
	wire [11:0] uncommitable_masks_2;

//AND all uncommittable mask
assign uncommitable_masks_2 = alu_T_2_uncom_2 &
div_r_uncom_2 & exe_reg_0_uncom_2 & exe_reg_1_uncom_2 & exe_reg_2_uncom_2 & rrd_0_uncom_2 &
rrd_1_uncom_2 & rrd_2_uncom_2 & bkq_0_uncom_2 & bkq_1_uncom_2 & bkq_2_uncom_2 &
bkq_3_uncom_2 & bkq_4_uncom_2 & alu_T_2_0_uncom_2 & alu_T_2_1_uncom_2 & alu_T_2_2_uncom_2 &
ifpu_T_2_0_uncom_2 & ifpu_T_2_1_uncom_2 & imul_T_2_0_uncom_2 & imul_T_2_1_uncom_2 &
imul_T_2_2_uncom_2 & fp_issue_slot_0_uncom_2 & fp_issue_slot_1_uncom_2 & fp_issue_slot_2_uncom_2 & fp_issue_slot_3_uncom_2 &
fp_issue_slot_4_uncom_2 & fp_issue_slot_5_uncom_2 & fp_issue_slot_6_uncom_2 & fp_issue_slot_7_uncom_2 & fp_issue_slot_8_uncom_2 &
fp_issue_slot_9_uncom_2 & fp_issue_slot_10_uncom_2 & fp_issue_slot_11_uncom_2 & fp_issue_slot_12_uncom_2 & fp_issue_slot_13_uncom_2 &
fp_issue_slot_14_uncom_2 & fp_issue_slot_15_uncom_2 & fp_bkq_0_uncom_2 & fp_bkq_1_uncom_2 & fp_bkq_2_uncom_2 &
fp_bkq_3_uncom_2 & fp_bkq_4_uncom_2 & fp_bkq_5_uncom_2 & fp_bkq_6_uncom_2 & fp_bkq_1_0_uncom_2 &
fp_bkq_1_1_uncom_2 & fp_bkq_1_2_uncom_2 & fdiv_buf_uncom_2 & fdiv_divsqrt_uncom_2 & fdiv_out_uncom_2 &
fpu_T_2_0_uncom_2 & fpu_T_2_1_uncom_2 & fpu_T_2_2_uncom_2 & fpu_T_2_3_uncom_2 & f_exe_reg_uncom_2 &
f_rrd_uncom_2 & int_issue_slot_0_uncom_2 & int_issue_slot_1_uncom_2 & int_issue_slot_2_uncom_2 & int_issue_slot_3_uncom_2 &
int_issue_slot_4_uncom_2 & int_issue_slot_5_uncom_2 & int_issue_slot_6_uncom_2 & int_issue_slot_7_uncom_2 & int_issue_slot_8_uncom_2 &
int_issue_slot_9_uncom_2 & int_issue_slot_10_uncom_2 & int_issue_slot_11_uncom_2 & int_issue_slot_12_uncom_2 & int_issue_slot_13_uncom_2 &
int_issue_slot_14_uncom_2 & int_issue_slot_15_uncom_2 & int_issue_slot_16_uncom_2 & int_issue_slot_17_uncom_2 & int_issue_slot_18_uncom_2 &
int_issue_slot_19_uncom_2 & mem_issue_slot_0_uncom_2 & mem_issue_slot_1_uncom_2 & mem_issue_slot_2_uncom_2 & mem_issue_slot_3_uncom_2 &
mem_issue_slot_4_uncom_2 & mem_issue_slot_5_uncom_2 & mem_issue_slot_6_uncom_2 & mem_issue_slot_7_uncom_2 & mem_issue_slot_8_uncom_2 &
mem_issue_slot_9_uncom_2 & mem_issue_slot_10_uncom_2 & mem_issue_slot_11_uncom_2 & lsu_ldq_0_uncom_2 & lsu_ldq_1_uncom_2 &
lsu_ldq_2_uncom_2 & lsu_ldq_3_uncom_2 & lsu_ldq_4_uncom_2 & lsu_ldq_5_uncom_2 & lsu_ldq_6_uncom_2 &
lsu_ldq_7_uncom_2 & lsu_ldq_8_uncom_2 & lsu_ldq_9_uncom_2 & lsu_ldq_10_uncom_2 & lsu_ldq_11_uncom_2 &
lsu_ldq_12_uncom_2 & lsu_ldq_13_uncom_2 & lsu_ldq_14_uncom_2 & lsu_ldq_15_uncom_2 & lsu_mem_uncom_2 &
lsu_mem_stq_uncom_2 & lsu_mem_retry_uncom_2 & lsu_mem_xcpt_uncom_2 & lsu_stdf_uncom_2 & lsu_mem_stdf_uncom_2 & lsu_stq_0_uncom_2 &
lsu_stq_1_uncom_2 & lsu_stq_2_uncom_2 & lsu_stq_3_uncom_2 & lsu_stq_4_uncom_2 & lsu_stq_5_uncom_2 &
lsu_stq_6_uncom_2 & lsu_stq_7_uncom_2 & lsu_stq_8_uncom_2 & lsu_stq_9_uncom_2 & lsu_stq_10_uncom_2 &
lsu_stq_11_uncom_2 & lsu_stq_12_uncom_2 & lsu_stq_13_uncom_2 & lsu_stq_14_uncom_2 & lsu_stq_15_uncom_2 &
rob__0_uncom_2 & rob__1_uncom_2 & rob__2_uncom_2 & rob__3_uncom_2 & rob__4_uncom_2 &
rob__5_uncom_2 & rob__6_uncom_2 & rob__7_uncom_2 & rob__8_uncom_2 & rob__9_uncom_2 &
rob__10_uncom_2 & rob__11_uncom_2 & rob__12_uncom_2 & rob__13_uncom_2 & rob__14_uncom_2 &
rob__15_uncom_2 & rob__16_uncom_2 & rob__17_uncom_2 & rob__18_uncom_2 & rob__19_uncom_2 &
rob__20_uncom_2 & rob__21_uncom_2 & rob__22_uncom_2 & rob__23_uncom_2 & rob__24_uncom_2 &
rob__25_uncom_2 & rob__26_uncom_2 & rob__27_uncom_2 & rob__28_uncom_2 & rob__29_uncom_2 &
rob__30_uncom_2 & rob__31_uncom_2 & rob_1_0_uncom_2 & rob_1_1_uncom_2 & rob_1_2_uncom_2 &
rob_1_3_uncom_2 & rob_1_4_uncom_2 & rob_1_5_uncom_2 & rob_1_6_uncom_2 & rob_1_7_uncom_2 &
rob_1_8_uncom_2 & rob_1_9_uncom_2 & rob_1_10_uncom_2 & rob_1_11_uncom_2 & rob_1_12_uncom_2 &
rob_1_13_uncom_2 & rob_1_14_uncom_2 & rob_1_15_uncom_2 & rob_1_16_uncom_2 & rob_1_17_uncom_2 &
rob_1_18_uncom_2 & rob_1_19_uncom_2 & rob_1_20_uncom_2 & rob_1_21_uncom_2 & rob_1_22_uncom_2 &
rob_1_23_uncom_2 & rob_1_24_uncom_2 & rob_1_25_uncom_2 & rob_1_26_uncom_2 & rob_1_27_uncom_2 &
rob_1_28_uncom_2 & rob_1_29_uncom_2 & rob_1_30_uncom_2 & rob_1_31_uncom_2 &
lsu_clr_bsy_brmask_0_uncom_2 &
respq_uops_0_ldq_uncom_2 & respq_uops_1_ldq_uncom_2 & respq_uops_2_ldq_uncom_2 & respq_uops_3_ldq_uncom_2 &
respq_uops_0_stq_uncom_2 & respq_uops_1_stq_uncom_2 & respq_uops_2_stq_uncom_2 & respq_uops_3_stq_uncom_2 &
mmios_0_ldq_uncom_2 & mmios_0_stq_uncom_2 &
mshrs_0_rpq_uops_0_ldq_uncom_2 & mshrs_0_rpq_uops_1_ldq_uncom_2 & mshrs_0_rpq_uops_2_ldq_uncom_2 & mshrs_0_rpq_uops_3_ldq_uncom_2 &
mshrs_0_rpq_uops_4_ldq_uncom_2 & mshrs_0_rpq_uops_5_ldq_uncom_2 & mshrs_0_rpq_uops_6_ldq_uncom_2 & mshrs_0_rpq_uops_7_ldq_uncom_2 &
mshrs_0_rpq_uops_8_ldq_uncom_2 & mshrs_0_rpq_uops_9_ldq_uncom_2 & mshrs_0_rpq_uops_10_ldq_uncom_2 & mshrs_0_rpq_uops_11_ldq_uncom_2 &
mshrs_0_rpq_uops_12_ldq_uncom_2 & mshrs_0_rpq_uops_13_ldq_uncom_2 & mshrs_0_rpq_uops_14_ldq_uncom_2 & mshrs_0_rpq_uops_15_ldq_uncom_2 &/*
mshrs_0_rpq_uops_0_stq_uncom_2 & mshrs_0_rpq_uops_1_stq_uncom_2 & mshrs_0_rpq_uops_2_stq_uncom_2 & mshrs_0_rpq_uops_3_stq_uncom_2 &
mshrs_0_rpq_uops_4_stq_uncom_2 & mshrs_0_rpq_uops_5_stq_uncom_2 & mshrs_0_rpq_uops_6_stq_uncom_2 & mshrs_0_rpq_uops_7_stq_uncom_2 &
mshrs_0_rpq_uops_8_stq_uncom_2 & mshrs_0_rpq_uops_9_stq_uncom_2 & mshrs_0_rpq_uops_10_stq_uncom_2 & mshrs_0_rpq_uops_11_stq_uncom_2 &
mshrs_0_rpq_uops_12_stq_uncom_2 & mshrs_0_rpq_uops_13_stq_uncom_2 & mshrs_0_rpq_uops_14_stq_uncom_2 & mshrs_0_rpq_uops_15_stq_uncom_2 &*/
mshrs_1_rpq_uops_0_ldq_uncom_2 & mshrs_1_rpq_uops_1_ldq_uncom_2 & mshrs_1_rpq_uops_2_ldq_uncom_2 & mshrs_1_rpq_uops_3_ldq_uncom_2 &
mshrs_1_rpq_uops_4_ldq_uncom_2 & mshrs_1_rpq_uops_5_ldq_uncom_2 & mshrs_1_rpq_uops_6_ldq_uncom_2 & mshrs_1_rpq_uops_7_ldq_uncom_2 &
mshrs_1_rpq_uops_8_ldq_uncom_2 & mshrs_1_rpq_uops_9_ldq_uncom_2 & mshrs_1_rpq_uops_10_ldq_uncom_2 & mshrs_1_rpq_uops_11_ldq_uncom_2 &
mshrs_1_rpq_uops_12_ldq_uncom_2 & mshrs_1_rpq_uops_13_ldq_uncom_2 & mshrs_1_rpq_uops_14_ldq_uncom_2 & mshrs_1_rpq_uops_15_ldq_uncom_2 &/*
mshrs_1_rpq_uops_0_stq_uncom_2 & mshrs_1_rpq_uops_1_stq_uncom_2 & mshrs_1_rpq_uops_2_stq_uncom_2 & mshrs_1_rpq_uops_3_stq_uncom_2 &
mshrs_1_rpq_uops_4_stq_uncom_2 & mshrs_1_rpq_uops_5_stq_uncom_2 & mshrs_1_rpq_uops_6_stq_uncom_2 & mshrs_1_rpq_uops_7_stq_uncom_2 &
mshrs_1_rpq_uops_8_stq_uncom_2 & mshrs_1_rpq_uops_9_stq_uncom_2 & mshrs_1_rpq_uops_10_stq_uncom_2 & mshrs_1_rpq_uops_11_stq_uncom_2 &
mshrs_1_rpq_uops_12_stq_uncom_2 & mshrs_1_rpq_uops_13_stq_uncom_2 & mshrs_1_rpq_uops_14_stq_uncom_2 & mshrs_1_rpq_uops_15_stq_uncom_2 &*/
lsu_r_xcpt_uncom_2 & dcache_s1_req_ldq_uncom_2 &/* dcache_s1_req_stq_uncom_2 &*/ dcache_s2_req_ldq_uncom_2 /*& dcache_s2_req_stq_uncom_2*/;

//OR all committable masks
assign commitable_masks_2 = root_br_mask | alu_T_2_com_2 |
div_r_com_2 | exe_reg_0_com_2 | exe_reg_1_com_2 | exe_reg_2_com_2 | rrd_0_com_2 |
rrd_1_com_2 | rrd_2_com_2 | bkq_0_com_2 | bkq_1_com_2 | bkq_2_com_2 |
bkq_3_com_2 | bkq_4_com_2 | alu_T_2_0_com_2 | alu_T_2_1_com_2 | alu_T_2_2_com_2 |
ifpu_T_2_0_com_2 | ifpu_T_2_1_com_2 | imul_T_2_0_com_2 | imul_T_2_1_com_2 |
imul_T_2_2_com_2 | fp_issue_slot_0_com_2 | fp_issue_slot_1_com_2 | fp_issue_slot_2_com_2 | fp_issue_slot_3_com_2 |
fp_issue_slot_4_com_2 | fp_issue_slot_5_com_2 | fp_issue_slot_6_com_2 | fp_issue_slot_7_com_2 | fp_issue_slot_8_com_2 |
fp_issue_slot_9_com_2 | fp_issue_slot_10_com_2 | fp_issue_slot_11_com_2 | fp_issue_slot_12_com_2 | fp_issue_slot_13_com_2 |
fp_issue_slot_14_com_2 | fp_issue_slot_15_com_2 | fp_bkq_0_com_2 | fp_bkq_1_com_2 | fp_bkq_2_com_2 |
fp_bkq_3_com_2 | fp_bkq_4_com_2 | fp_bkq_5_com_2 | fp_bkq_6_com_2 | fp_bkq_1_0_com_2 |
fp_bkq_1_1_com_2 | fp_bkq_1_2_com_2 | fdiv_buf_com_2 | fdiv_divsqrt_com_2 | fdiv_out_com_2 |
fpu_T_2_0_com_2 | fpu_T_2_1_com_2 | fpu_T_2_2_com_2 | fpu_T_2_3_com_2 | f_exe_reg_com_2 |
f_rrd_com_2 | int_issue_slot_0_com_2 | int_issue_slot_1_com_2 | int_issue_slot_2_com_2 | int_issue_slot_3_com_2 |
int_issue_slot_4_com_2 | int_issue_slot_5_com_2 | int_issue_slot_6_com_2 | int_issue_slot_7_com_2 | int_issue_slot_8_com_2 |
int_issue_slot_9_com_2 | int_issue_slot_10_com_2 | int_issue_slot_11_com_2 | int_issue_slot_12_com_2 | int_issue_slot_13_com_2 |
int_issue_slot_14_com_2 | int_issue_slot_15_com_2 | int_issue_slot_16_com_2 | int_issue_slot_17_com_2 | int_issue_slot_18_com_2 |
int_issue_slot_19_com_2 | mem_issue_slot_0_com_2 | mem_issue_slot_1_com_2 | mem_issue_slot_2_com_2 | mem_issue_slot_3_com_2 |
mem_issue_slot_4_com_2 | mem_issue_slot_5_com_2 | mem_issue_slot_6_com_2 | mem_issue_slot_7_com_2 | mem_issue_slot_8_com_2 |
mem_issue_slot_9_com_2 | mem_issue_slot_10_com_2 | mem_issue_slot_11_com_2 | lsu_ldq_0_com_2 | lsu_ldq_1_com_2 |
lsu_ldq_2_com_2 | lsu_ldq_3_com_2 | lsu_ldq_4_com_2 | lsu_ldq_5_com_2 | lsu_ldq_6_com_2 |
lsu_ldq_7_com_2 | lsu_ldq_8_com_2 | lsu_ldq_9_com_2 | lsu_ldq_10_com_2 | lsu_ldq_11_com_2 |
lsu_ldq_12_com_2 | lsu_ldq_13_com_2 | lsu_ldq_14_com_2 | lsu_ldq_15_com_2 | lsu_mem_com_2 |
lsu_mem_stq_com_2 | lsu_mem_retry_com_2 | lsu_mem_xcpt_com_2 | lsu_stdf_com_2 | lsu_mem_stdf_com_2 | lsu_stq_0_com_2 |
lsu_stq_1_com_2 | lsu_stq_2_com_2 | lsu_stq_3_com_2 | lsu_stq_4_com_2 | lsu_stq_5_com_2 |
lsu_stq_6_com_2 | lsu_stq_7_com_2 | lsu_stq_8_com_2 | lsu_stq_9_com_2 | lsu_stq_10_com_2 |
lsu_stq_11_com_2 | lsu_stq_12_com_2 | lsu_stq_13_com_2 | lsu_stq_14_com_2 | lsu_stq_15_com_2 |
rob__0_com_2 | rob__1_com_2 | rob__2_com_2 | rob__3_com_2 | rob__4_com_2 |
rob__5_com_2 | rob__6_com_2 | rob__7_com_2 | rob__8_com_2 | rob__9_com_2 |
rob__10_com_2 | rob__11_com_2 | rob__12_com_2 | rob__13_com_2 | rob__14_com_2 |
rob__15_com_2 | rob__16_com_2 | rob__17_com_2 | rob__18_com_2 | rob__19_com_2 |
rob__20_com_2 | rob__21_com_2 | rob__22_com_2 | rob__23_com_2 | rob__24_com_2 |
rob__25_com_2 | rob__26_com_2 | rob__27_com_2 | rob__28_com_2 | rob__29_com_2 |
rob__30_com_2 | rob__31_com_2 | rob_1_0_com_2 | rob_1_1_com_2 | rob_1_2_com_2 |
rob_1_3_com_2 | rob_1_4_com_2 | rob_1_5_com_2 | rob_1_6_com_2 | rob_1_7_com_2 |
rob_1_8_com_2 | rob_1_9_com_2 | rob_1_10_com_2 | rob_1_11_com_2 | rob_1_12_com_2 |
rob_1_13_com_2 | rob_1_14_com_2 | rob_1_15_com_2 | rob_1_16_com_2 | rob_1_17_com_2 |
rob_1_18_com_2 | rob_1_19_com_2 | rob_1_20_com_2 | rob_1_21_com_2 | rob_1_22_com_2 |
rob_1_23_com_2 | rob_1_24_com_2 | rob_1_25_com_2 | rob_1_26_com_2 | rob_1_27_com_2 |
rob_1_28_com_2 | rob_1_29_com_2 | rob_1_30_com_2 | rob_1_31_com_2 |
lsu_clr_bsy_brmask_0_com_2 |
respq_uops_0_ldq_com_2 | respq_uops_1_ldq_com_2 | respq_uops_2_ldq_com_2 | respq_uops_3_ldq_com_2 |
respq_uops_0_stq_com_2 | respq_uops_1_stq_com_2 | respq_uops_2_stq_com_2 | respq_uops_3_stq_com_2 |
mmios_0_ldq_com_2 | mmios_0_stq_com_2 |
mshrs_0_rpq_uops_0_ldq_com_2 | mshrs_0_rpq_uops_1_ldq_com_2 | mshrs_0_rpq_uops_2_ldq_com_2 | mshrs_0_rpq_uops_3_ldq_com_2 |
mshrs_0_rpq_uops_4_ldq_com_2 | mshrs_0_rpq_uops_5_ldq_com_2 | mshrs_0_rpq_uops_6_ldq_com_2 | mshrs_0_rpq_uops_7_ldq_com_2 |
mshrs_0_rpq_uops_8_ldq_com_2 | mshrs_0_rpq_uops_9_ldq_com_2 | mshrs_0_rpq_uops_10_ldq_com_2 | mshrs_0_rpq_uops_11_ldq_com_2 |
mshrs_0_rpq_uops_12_ldq_com_2 | mshrs_0_rpq_uops_13_ldq_com_2 | mshrs_0_rpq_uops_14_ldq_com_2 | mshrs_0_rpq_uops_15_ldq_com_2 |/*
mshrs_0_rpq_uops_0_stq_com_2 | mshrs_0_rpq_uops_1_stq_com_2 | mshrs_0_rpq_uops_2_stq_com_2 | mshrs_0_rpq_uops_3_stq_com_2 |
mshrs_0_rpq_uops_4_stq_com_2 | mshrs_0_rpq_uops_5_stq_com_2 | mshrs_0_rpq_uops_6_stq_com_2 | mshrs_0_rpq_uops_7_stq_com_2 |
mshrs_0_rpq_uops_8_stq_com_2 | mshrs_0_rpq_uops_9_stq_com_2 | mshrs_0_rpq_uops_10_stq_com_2 | mshrs_0_rpq_uops_11_stq_com_2 |
mshrs_0_rpq_uops_12_stq_com_2 | mshrs_0_rpq_uops_13_stq_com_2 | mshrs_0_rpq_uops_14_stq_com_2 | mshrs_0_rpq_uops_15_stq_com_2 |*/
mshrs_1_rpq_uops_0_ldq_com_2 | mshrs_1_rpq_uops_1_ldq_com_2 | mshrs_1_rpq_uops_2_ldq_com_2 | mshrs_1_rpq_uops_3_ldq_com_2 |
mshrs_1_rpq_uops_4_ldq_com_2 | mshrs_1_rpq_uops_5_ldq_com_2 | mshrs_1_rpq_uops_6_ldq_com_2 | mshrs_1_rpq_uops_7_ldq_com_2 |
mshrs_1_rpq_uops_8_ldq_com_2 | mshrs_1_rpq_uops_9_ldq_com_2 | mshrs_1_rpq_uops_10_ldq_com_2 | mshrs_1_rpq_uops_11_ldq_com_2 |
mshrs_1_rpq_uops_12_ldq_com_2 | mshrs_1_rpq_uops_13_ldq_com_2 | mshrs_1_rpq_uops_14_ldq_com_2 | mshrs_1_rpq_uops_15_ldq_com_2 |/*
mshrs_1_rpq_uops_0_stq_com_2 | mshrs_1_rpq_uops_1_stq_com_2 | mshrs_1_rpq_uops_2_stq_com_2 | mshrs_1_rpq_uops_3_stq_com_2 |
mshrs_1_rpq_uops_4_stq_com_2 | mshrs_1_rpq_uops_5_stq_com_2 | mshrs_1_rpq_uops_6_stq_com_2 | mshrs_1_rpq_uops_7_stq_com_2 |
mshrs_1_rpq_uops_8_stq_com_2 | mshrs_1_rpq_uops_9_stq_com_2 | mshrs_1_rpq_uops_10_stq_com_2 | mshrs_1_rpq_uops_11_stq_com_2 |
mshrs_1_rpq_uops_12_stq_com_2 | mshrs_1_rpq_uops_13_stq_com_2 | mshrs_1_rpq_uops_14_stq_com_2 | mshrs_1_rpq_uops_15_stq_com_2 |*/
lsu_r_xcpt_com_2 | dcache_s1_req_ldq_com_2 | /*dcache_s1_req_stq_com_2 |*/ dcache_s2_req_ldq_com_2 /*| dcache_s2_req_stq_com_2*/;

//****************************************************//
//************ME-5(Consistent Speculation Tag)********//

	wire [11:0] uncommitable_masks;
	wire ME_5;

  //combine uncommittable masks of both SoCs
	assign uncommitable_masks = uncommitable_masks_1 & uncommitable_masks_2;

  //all uncommittable masks must have the same bit set as root_br_mask
  //this means that every uncommittable instruction is speculated under the instruction at root_ID
	assign ME_5 = ( ((mispred_happened_1 == 1'b1) && (mispred_happened_2 == 1'b1)) || root_id_killed || root_id_already_killed || (uncommitable_masks & root_br_mask) == root_br_mask );

//****************************************************//
//************ME-6(Consistent Spawn Tag)**************//


	wire ME_6_1;
	wire ME_6_2;
	wire ME_6;

	//if a branch is resolved, its ROB ID must either be in the committable set or it must have a spawn tag greater than T_main
  //changed to: check for all buffers if the contained branch is either in the committable set or has a spawn tag greater than T_main
	assign ME_6_1 = ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed))
                  ?
                  (
                  ((soc1.core.b2_mispredict == 1'b1) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.b2_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.b2_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.brinfos_0_valid == 1'b1) && (soc1.core.brinfos_0_mispredict == 1'b1) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.brinfos_0_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.brinfos_0_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.brinfos_1_valid == 1'b1) && (soc1.core.brinfos_1_mispredict == 1'b1) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.brinfos_1_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.brinfos_1_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_0.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_0.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_0.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_1.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_1.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_1.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_2.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_2.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_2.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_3.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_3.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_3.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_4.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_4.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_4.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_5.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_5.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_5.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_6.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_6.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_6.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_7.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_7.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_7.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_8.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_8.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_8.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_9.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_9.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_9.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_10.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_10.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_10.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_11.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_11.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_11.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_12.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_12.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_12.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_13.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_13.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_13.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_14.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_14.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_14.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_15.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_15.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_15.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_16.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_16.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_16.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_17.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_17.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_17.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_18.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_18.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_18.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.int_issue_unit.slots_19.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.int_issue_unit.slots_19.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.int_issue_unit.slots_19.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  (soc1.core.iregister_read.exe_reg_valids_1 && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.exe_reg_uops_1_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.iregister_read.exe_reg_uops_1_br_tag, commitable_masks_1) : 1'b1) &&
                  (soc1.core.iregister_read.exe_reg_valids_2 && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.exe_reg_uops_2_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.iregister_read.exe_reg_uops_2_br_tag, commitable_masks_1) : 1'b1) &&
                  (soc1.core.iregister_read.rrd_valids_1_REG && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.rrd_uops_1_REG_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.iregister_read.rrd_uops_1_REG_br_tag, commitable_masks_1) : 1'b1) &&
                  (soc1.core.iregister_read.rrd_valids_2_REG && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.iregister_read.rrd_uops_2_REG_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.iregister_read.rrd_uops_2_REG_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_0.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_0.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_0.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_1.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_1.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_1.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_2.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_2.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_2.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_3.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_3.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_3.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_4.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_4.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_4.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_5.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_5.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_5.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_6.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_6.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_6.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_7.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_7.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_7.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_8.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_8.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_8.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_9.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_9.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_9.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_10.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_10.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_10.slot_uop_br_tag, commitable_masks_1) : 1'b1) &&
                  ((soc1.core.mem_issue_unit.slots_11.state != 2'b0) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.mem_issue_unit.slots_11.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc1.core.mem_issue_unit.slots_11.slot_uop_br_tag, commitable_masks_1) : 1'b1))
                  :
                  1'b1
                  ;

	assign ME_6_2 = ((mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) && (!root_id_killed && !root_id_already_killed))
                  ?
                  (
                  ((soc2.core.b2_mispredict == 1'b1) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.b2_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.b2_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.brinfos_0_valid == 1'b1) && (soc2.core.brinfos_0_mispredict == 1'b1) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.brinfos_0_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.brinfos_0_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.brinfos_1_valid == 1'b1) && (soc2.core.brinfos_1_mispredict == 1'b1) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.brinfos_1_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.brinfos_1_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_0.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_0.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_0.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_1.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_1.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_1.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_2.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_2.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_2.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_3.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_3.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_3.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_4.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_4.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_4.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_5.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_5.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_5.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_6.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_6.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_6.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_7.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_7.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_7.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_8.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_8.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_8.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_9.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_9.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_9.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_10.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_10.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_10.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_11.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_11.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_11.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_12.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_12.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_12.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_13.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_13.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_13.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_14.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_14.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_14.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_15.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_15.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_15.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_16.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_16.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_16.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_17.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_17.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_17.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_18.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_18.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_18.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.int_issue_unit.slots_19.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.int_issue_unit.slots_19.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.int_issue_unit.slots_19.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  (soc2.core.iregister_read.exe_reg_valids_1 && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.exe_reg_uops_1_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.iregister_read.exe_reg_uops_1_br_tag, commitable_masks_2) : 1'b1) &&
                  (soc2.core.iregister_read.exe_reg_valids_2 && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.exe_reg_uops_2_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.iregister_read.exe_reg_uops_2_br_tag, commitable_masks_2) : 1'b1) &&
                  (soc2.core.iregister_read.rrd_valids_1_REG && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.rrd_uops_1_REG_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.iregister_read.rrd_uops_1_REG_br_tag, commitable_masks_2) : 1'b1) &&
                  (soc2.core.iregister_read.rrd_valids_2_REG && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.iregister_read.rrd_uops_2_REG_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.iregister_read.rrd_uops_2_REG_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_0.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_0.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_0.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_1.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_1.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_1.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_2.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_2.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_2.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_3.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_3.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_3.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_4.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_4.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_4.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_5.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_5.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_5.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_6.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_6.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_6.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_7.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_7.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_7.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_8.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_8.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_8.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_9.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_9.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_9.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_10.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_10.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_10.slot_uop_br_tag, commitable_masks_2) : 1'b1) &&
                  ((soc2.core.mem_issue_unit.slots_11.state != 2'b0) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.mem_issue_unit.slots_11.slot_uop_rob_idx) != 1'b1) ?
                      isSpawnTagGreater(soc2.core.mem_issue_unit.slots_11.slot_uop_br_tag, commitable_masks_2) : 1'b1))
                  :
                  1'b1
                  ;

	assign ME_6 = ME_6_1 && ME_6_2;

//****************************************************//
//************MicroEquivalence************************//

	wire microequivalence;

	assign microequivalence = ME_1 && ME_2 && ME_3 && ME_4 && ME_5 && ME_6;

//****************************************************//
//************L-Alert Definition**********************//

  wire root_id_killed;
  assign root_id_killed =
  !(
    ((soc1.core.rob.rob_head < soc1.core.rob.rob_tail) && (soc1.core.rob.rob_head <= root_id[5:1]) && (root_id[5:1] < soc1.core.rob.rob_tail)||
    !(soc1.core.rob.rob_head < soc1.core.rob.rob_tail) && (soc1.core.rob.rob_head > soc1.core.rob.rob_tail) && ((soc1.core.rob.rob_head <= root_id[5:1]) || (root_id[5:1] < soc1.core.rob.rob_tail))||
    !(soc1.core.rob.rob_head < soc1.core.rob.rob_tail) && !(soc1.core.rob.rob_head > soc1.core.rob.rob_tail) && !soc1.core.rob.io_empty) &&
    rob_valids_1[root_id]
   ) &&

  !(
    ((soc2.core.rob.rob_head < soc2.core.rob.rob_tail) && (soc2.core.rob.rob_head <= root_id[5:1]) && (root_id[5:1] < soc2.core.rob.rob_tail)||
    !(soc2.core.rob.rob_head < soc2.core.rob.rob_tail) && (soc2.core.rob.rob_head > soc2.core.rob.rob_tail) && ((soc2.core.rob.rob_head <= root_id[5:1]) || (root_id[5:1] < soc2.core.rob.rob_tail))||
    !(soc2.core.rob.rob_head < soc2.core.rob.rob_tail) && !(soc2.core.rob.rob_head > soc2.core.rob.rob_tail) && !soc2.core.rob.io_empty) &&
    rob_valids_2[root_id]
   );

  reg root_id_already_killed;

  always @(posedge clock)
    begin
      if (reset)
      begin
        root_id_already_killed <= 1'b0;
      end
      else
      begin
        if(root_id_killed == 1'b1)
        begin
          root_id_already_killed <= 1'b1;
        end
      end
    end

	wire lAlert;

	assign lAlert = !(mispred_happened_1 && mispred_happened_2) && (!root_id_killed && !root_id_already_killed) && (soc1.core.rob.io_commit_valids_0 != soc2.core.rob.io_commit_valids_0 || soc1.core.rob.io_commit_valids_1 != soc2.core.rob.io_commit_valids_1);

	wire lAlert_earlyAlarm;
	assign lAlert_earlyAlarm = mispred_flag_1 != mispred_flag_2;
	
	wire pnr_between_head_and_root_id;
	assign pnr_between_head_and_root_id = 
		!(mispred_happened_1 && mispred_happened_2) && (!root_id_killed && !root_id_already_killed)
		?
			ROBisOlder(soc1.core.rob.io_rob_pnr_idx, root_id, soc1.core.rob.io_rob_head_idx) || (soc1.core.rob.io_rob_pnr_idx == root_id) &&
			ROBisOlder(soc2.core.rob.io_rob_pnr_idx, root_id, soc2.core.rob.io_rob_head_idx) || (soc2.core.rob.io_rob_pnr_idx == root_id)
		:
			1'b1;
	;
	
	wire tainted_lsu_resp_rob_idx_and_yrot_equal;
	assign tainted_lsu_resp_rob_idx_and_yrot_equal = 
		(soc1.lsu.io_core_exe_0_iresp_bits_uop_taint && soc1.lsu.io_core_exe_0_iresp_valid ? soc1.lsu.io_core_exe_0_iresp_bits_uop_rob_idx == soc1.lsu.io_core_exe_0_iresp_bits_uop_yrot : 1'b1) &&
		(soc2.lsu.io_core_exe_0_iresp_bits_uop_taint && soc2.lsu.io_core_exe_0_iresp_valid ? soc2.lsu.io_core_exe_0_iresp_bits_uop_rob_idx == soc2.lsu.io_core_exe_0_iresp_bits_uop_yrot : 1'b1) &&
		(soc1.lsu.io_core_exe_0_fresp_bits_uop_taint && soc1.lsu.io_core_exe_0_fresp_valid ? soc1.lsu.io_core_exe_0_fresp_bits_uop_rob_idx == soc1.lsu.io_core_exe_0_fresp_bits_uop_yrot : 1'b1) &&
		(soc2.lsu.io_core_exe_0_fresp_bits_uop_taint && soc2.lsu.io_core_exe_0_fresp_valid ? soc2.lsu.io_core_exe_0_fresp_bits_uop_rob_idx == soc2.lsu.io_core_exe_0_fresp_bits_uop_yrot : 1'b1)
	;
	

  //recursive definition of committable elements relative to head
  //an element is committable if its rob_idx is committable and all prior elements until head are committable
  wire is_stq1_committable_head_0;
  assign is_stq1_committable_head_0 = isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[soc1.lsu.stq_head]);
  wire is_stq1_committable_head_1;
  assign is_stq1_committable_head_1 = is_stq1_committable_head_0 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +1) % 16]);
  wire is_stq1_committable_head_2;
  assign is_stq1_committable_head_2 = is_stq1_committable_head_1 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +2) % 16]);
  wire is_stq1_committable_head_3;
  assign is_stq1_committable_head_3 = is_stq1_committable_head_2 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +3) % 16]);
  wire is_stq1_committable_head_4;
  assign is_stq1_committable_head_4 = is_stq1_committable_head_3 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +4) % 16]);
  wire is_stq1_committable_head_5;
  assign is_stq1_committable_head_5 = is_stq1_committable_head_4 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +5) % 16]);
  wire is_stq1_committable_head_6;
  assign is_stq1_committable_head_6 = is_stq1_committable_head_5 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +6) % 16]);
  wire is_stq1_committable_head_7;
  assign is_stq1_committable_head_7 = is_stq1_committable_head_6 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +7) % 16]);
  wire is_stq1_committable_head_8;
  assign is_stq1_committable_head_8 = is_stq1_committable_head_7 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +8) % 16]);
  wire is_stq1_committable_head_9;
  assign is_stq1_committable_head_9 = is_stq1_committable_head_8 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +9) % 16]);
  wire is_stq1_committable_head_10;
  assign is_stq1_committable_head_10 = is_stq1_committable_head_9 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +10) % 16]);
  wire is_stq1_committable_head_11;
  assign is_stq1_committable_head_11 = is_stq1_committable_head_10 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +11) % 16]);
  wire is_stq1_committable_head_12;
  assign is_stq1_committable_head_12 = is_stq1_committable_head_11 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +12) % 16]);
  wire is_stq1_committable_head_13;
  assign is_stq1_committable_head_13 = is_stq1_committable_head_12 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +13) % 16]);
  wire is_stq1_committable_head_14;
  assign is_stq1_committable_head_14 = is_stq1_committable_head_13 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +14) % 16]);
  wire is_stq1_committable_head_15;
  assign is_stq1_committable_head_15 = is_stq1_committable_head_14 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, stq_rob_idx_1[(soc1.lsu.stq_head +15) % 16]);

  //recursive definition of committable elements relative to head
  //an element is committable if its rob_idx is committable and all prior elements until head are committable
  wire is_stq2_committable_head_0;
  assign is_stq2_committable_head_0 = isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[soc2.lsu.stq_head]);
  wire is_stq2_committable_head_1;
  assign is_stq2_committable_head_1 = is_stq2_committable_head_0 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +1) % 16]);
  wire is_stq2_committable_head_2;
  assign is_stq2_committable_head_2 = is_stq2_committable_head_1 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +2) % 16]);
  wire is_stq2_committable_head_3;
  assign is_stq2_committable_head_3 = is_stq2_committable_head_2 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +3) % 16]);
  wire is_stq2_committable_head_4;
  assign is_stq2_committable_head_4 = is_stq2_committable_head_3 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +4) % 16]);
  wire is_stq2_committable_head_5;
  assign is_stq2_committable_head_5 = is_stq2_committable_head_4 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +5) % 16]);
  wire is_stq2_committable_head_6;
  assign is_stq2_committable_head_6 = is_stq2_committable_head_5 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +6) % 16]);
  wire is_stq2_committable_head_7;
  assign is_stq2_committable_head_7 = is_stq2_committable_head_6 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +7) % 16]);
  wire is_stq2_committable_head_8;
  assign is_stq2_committable_head_8 = is_stq2_committable_head_7 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +8) % 16]);
  wire is_stq2_committable_head_9;
  assign is_stq2_committable_head_9 = is_stq2_committable_head_8 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +9) % 16]);
  wire is_stq2_committable_head_10;
  assign is_stq2_committable_head_10 = is_stq2_committable_head_9 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +10) % 16]);
  wire is_stq2_committable_head_11;
  assign is_stq2_committable_head_11 = is_stq2_committable_head_10 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +11) % 16]);
  wire is_stq2_committable_head_12;
  assign is_stq2_committable_head_12 = is_stq2_committable_head_11 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +12) % 16]);
  wire is_stq2_committable_head_13;
  assign is_stq2_committable_head_13 = is_stq2_committable_head_12 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +13) % 16]);
  wire is_stq2_committable_head_14;
  assign is_stq2_committable_head_14 = is_stq2_committable_head_13 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +14) % 16]);
  wire is_stq2_committable_head_15;
  assign is_stq2_committable_head_15 = is_stq2_committable_head_14 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, stq_rob_idx_2[(soc2.lsu.stq_head +15) % 16]);

  //function that maps the rob_idx to the "head-relative" entry
  function automatic is_stq1_committable;
    //4-bit ID of the store queue entry
    input [3:0] idx;
    begin
      //mapping: (position of entry relative to head) -> (actual index of entry)
      case(idx)
        soc1.lsu.stq_head         : is_stq1_committable = is_stq1_committable_head_0;
        (soc1.lsu.stq_head+1)%16  : is_stq1_committable = is_stq1_committable_head_1;
        (soc1.lsu.stq_head+2)%16  : is_stq1_committable = is_stq1_committable_head_2;
        (soc1.lsu.stq_head+3)%16  : is_stq1_committable = is_stq1_committable_head_3;
        (soc1.lsu.stq_head+4)%16  : is_stq1_committable = is_stq1_committable_head_4;
        (soc1.lsu.stq_head+5)%16  : is_stq1_committable = is_stq1_committable_head_5;
        (soc1.lsu.stq_head+6)%16  : is_stq1_committable = is_stq1_committable_head_6;
        (soc1.lsu.stq_head+7)%16  : is_stq1_committable = is_stq1_committable_head_7;
        (soc1.lsu.stq_head+8)%16  : is_stq1_committable = is_stq1_committable_head_8;
        (soc1.lsu.stq_head+9)%16  : is_stq1_committable = is_stq1_committable_head_9;
        (soc1.lsu.stq_head+10)%16 : is_stq1_committable = is_stq1_committable_head_10;
        (soc1.lsu.stq_head+11)%16 : is_stq1_committable = is_stq1_committable_head_11;
        (soc1.lsu.stq_head+12)%16 : is_stq1_committable = is_stq1_committable_head_12;
        (soc1.lsu.stq_head+13)%16 : is_stq1_committable = is_stq1_committable_head_13;
        (soc1.lsu.stq_head+14)%16 : is_stq1_committable = is_stq1_committable_head_14;
        (soc1.lsu.stq_head+15)%16 : is_stq1_committable = is_stq1_committable_head_15;
        default                   : is_stq1_committable = 1'b0;
      endcase
    end
  endfunction

  //function that maps the rob_idx to the "head-relative" entry
  function automatic is_stq2_committable;
    //4-bit ID of the store queue entry
    input [3:0] idx;
    begin
      //mapping: (position of entry relative to head) -> (actual index of entry)
      case(idx)
        soc2.lsu.stq_head         : is_stq2_committable = is_stq2_committable_head_0;
        (soc2.lsu.stq_head+1)%16  : is_stq2_committable = is_stq2_committable_head_1;
        (soc2.lsu.stq_head+2)%16  : is_stq2_committable = is_stq2_committable_head_2;
        (soc2.lsu.stq_head+3)%16  : is_stq2_committable = is_stq2_committable_head_3;
        (soc2.lsu.stq_head+4)%16  : is_stq2_committable = is_stq2_committable_head_4;
        (soc2.lsu.stq_head+5)%16  : is_stq2_committable = is_stq2_committable_head_5;
        (soc2.lsu.stq_head+6)%16  : is_stq2_committable = is_stq2_committable_head_6;
        (soc2.lsu.stq_head+7)%16  : is_stq2_committable = is_stq2_committable_head_7;
        (soc2.lsu.stq_head+8)%16  : is_stq2_committable = is_stq2_committable_head_8;
        (soc2.lsu.stq_head+9)%16  : is_stq2_committable = is_stq2_committable_head_9;
        (soc2.lsu.stq_head+10)%16 : is_stq2_committable = is_stq2_committable_head_10;
        (soc2.lsu.stq_head+11)%16 : is_stq2_committable = is_stq2_committable_head_11;
        (soc2.lsu.stq_head+12)%16 : is_stq2_committable = is_stq2_committable_head_12;
        (soc2.lsu.stq_head+13)%16 : is_stq2_committable = is_stq2_committable_head_13;
        (soc2.lsu.stq_head+14)%16 : is_stq2_committable = is_stq2_committable_head_14;
        (soc2.lsu.stq_head+15)%16 : is_stq2_committable = is_stq2_committable_head_15;
        default                   : is_stq2_committable = 1'b0;
      endcase
    end
  endfunction

	wire [15:0] stq1_0_st_dep_mask;
	wire [15:0] stq1_1_st_dep_mask;
	wire [15:0] stq1_2_st_dep_mask;
	wire [15:0] stq1_3_st_dep_mask;
	wire [15:0] stq1_4_st_dep_mask;
	wire [15:0] stq1_5_st_dep_mask;
	wire [15:0] stq1_6_st_dep_mask;
	wire [15:0] stq1_7_st_dep_mask;
	wire [15:0] stq1_8_st_dep_mask;
	wire [15:0] stq1_9_st_dep_mask;
	wire [15:0] stq1_10_st_dep_mask;
	wire [15:0] stq1_11_st_dep_mask;
	wire [15:0] stq1_12_st_dep_mask;
	wire [15:0] stq1_13_st_dep_mask;
	wire [15:0] stq1_14_st_dep_mask;
	wire [15:0] stq1_15_st_dep_mask;

  //create the dependency masks for all stores that are uncommittable
	assign stq1_0_st_dep_mask = is_stq1_committable(4'b0000) ? 16'b0 : (16'b1 << 0);
	assign stq1_1_st_dep_mask = is_stq1_committable(4'b0001) ? 16'b0 : (16'b1 << 1);
	assign stq1_2_st_dep_mask = is_stq1_committable(4'b0010) ? 16'b0 : (16'b1 << 2);
	assign stq1_3_st_dep_mask = is_stq1_committable(4'b0011) ? 16'b0 : (16'b1 << 3);
	assign stq1_4_st_dep_mask = is_stq1_committable(4'b0100) ? 16'b0 : (16'b1 << 4);
	assign stq1_5_st_dep_mask = is_stq1_committable(4'b0101) ? 16'b0 : (16'b1 << 5);
	assign stq1_6_st_dep_mask = is_stq1_committable(4'b0110) ? 16'b0 : (16'b1 << 6);
	assign stq1_7_st_dep_mask = is_stq1_committable(4'b0111) ? 16'b0 : (16'b1 << 7);
	assign stq1_8_st_dep_mask = is_stq1_committable(4'b1000) ? 16'b0 : (16'b1 << 8);
	assign stq1_9_st_dep_mask = is_stq1_committable(4'b1001) ? 16'b0 : (16'b1 << 9);
	assign stq1_10_st_dep_mask = is_stq1_committable(4'b1010) ? 16'b0 : (16'b1 << 10);
	assign stq1_11_st_dep_mask = is_stq1_committable(4'b1011) ? 16'b0 : (16'b1 << 11);
	assign stq1_12_st_dep_mask = is_stq1_committable(4'b1100) ? 16'b0 : (16'b1 << 12);
	assign stq1_13_st_dep_mask = is_stq1_committable(4'b1101) ? 16'b0 : (16'b1 << 13);
	assign stq1_14_st_dep_mask = is_stq1_committable(4'b1110) ? 16'b0 : (16'b1 << 14);
	assign stq1_15_st_dep_mask = is_stq1_committable(4'b1111) ? 16'b0 : (16'b1 << 15);

  //OR the st_dep_masks of all uncommittable stores
	wire [15:0] uncom1_st_dep_mask;
	assign uncom1_st_dep_mask = stq1_0_st_dep_mask | stq1_1_st_dep_mask | stq1_2_st_dep_mask | stq1_3_st_dep_mask |
	stq1_4_st_dep_mask | stq1_5_st_dep_mask | stq1_6_st_dep_mask | stq1_7_st_dep_mask | stq1_8_st_dep_mask |
	stq1_9_st_dep_mask | stq1_10_st_dep_mask | stq1_11_st_dep_mask | stq1_12_st_dep_mask | stq1_13_st_dep_mask | stq1_14_st_dep_mask | stq1_15_st_dep_mask;

  wire [15:0] stq2_0_st_dep_mask;
	wire [15:0] stq2_1_st_dep_mask;
	wire [15:0] stq2_2_st_dep_mask;
	wire [15:0] stq2_3_st_dep_mask;
	wire [15:0] stq2_4_st_dep_mask;
	wire [15:0] stq2_5_st_dep_mask;
	wire [15:0] stq2_6_st_dep_mask;
	wire [15:0] stq2_7_st_dep_mask;
	wire [15:0] stq2_8_st_dep_mask;
	wire [15:0] stq2_9_st_dep_mask;
	wire [15:0] stq2_10_st_dep_mask;
	wire [15:0] stq2_11_st_dep_mask;
	wire [15:0] stq2_12_st_dep_mask;
	wire [15:0] stq2_13_st_dep_mask;
	wire [15:0] stq2_14_st_dep_mask;
	wire [15:0] stq2_15_st_dep_mask;

  //create the dependency masks for all stores that are uncommittable
	assign stq2_0_st_dep_mask = is_stq2_committable(4'b0000) ? 16'b0 : 16'b1 << 0;
	assign stq2_1_st_dep_mask = is_stq2_committable(4'b0001) ? 16'b0 : 16'b1 << 1;
	assign stq2_2_st_dep_mask = is_stq2_committable(4'b0010) ? 16'b0 : 16'b1 << 2;
	assign stq2_3_st_dep_mask = is_stq2_committable(4'b0011) ? 16'b0 : 16'b1 << 3;
	assign stq2_4_st_dep_mask = is_stq2_committable(4'b0100) ? 16'b0 : 16'b1 << 4;
	assign stq2_5_st_dep_mask = is_stq2_committable(4'b0101) ? 16'b0 : 16'b1 << 5;
	assign stq2_6_st_dep_mask = is_stq2_committable(4'b0110) ? 16'b0 : 16'b1 << 6;
	assign stq2_7_st_dep_mask = is_stq2_committable(4'b0111) ? 16'b0 : 16'b1 << 7;
	assign stq2_8_st_dep_mask = is_stq2_committable(4'b1000) ? 16'b0 : 16'b1 << 8;
	assign stq2_9_st_dep_mask = is_stq2_committable(4'b1001) ? 16'b0 : 16'b1 << 9;
	assign stq2_10_st_dep_mask = is_stq2_committable(4'b1010) ? 16'b0 : 16'b1 << 10;
	assign stq2_11_st_dep_mask = is_stq2_committable(4'b1011) ? 16'b0 : 16'b1 << 11;
	assign stq2_12_st_dep_mask = is_stq2_committable(4'b1100) ? 16'b0 : 16'b1 << 12;
	assign stq2_13_st_dep_mask = is_stq2_committable(4'b1101) ? 16'b0 : 16'b1 << 13;
	assign stq2_14_st_dep_mask = is_stq2_committable(4'b1110) ? 16'b0 : 16'b1 << 14;
	assign stq2_15_st_dep_mask = is_stq2_committable(4'b1111) ? 16'b0 : 16'b1 << 15;

  //OR the st_dep_masks of all uncommittable stores
	wire [15:0] uncom2_st_dep_mask;
	assign uncom2_st_dep_mask = stq2_0_st_dep_mask | stq2_1_st_dep_mask | stq2_2_st_dep_mask | stq2_3_st_dep_mask |
	stq2_4_st_dep_mask | stq2_5_st_dep_mask | stq2_6_st_dep_mask | stq2_7_st_dep_mask | stq2_8_st_dep_mask |
	stq2_9_st_dep_mask | stq2_10_st_dep_mask | stq2_11_st_dep_mask | stq2_12_st_dep_mask | stq2_13_st_dep_mask | stq2_14_st_dep_mask | stq2_15_st_dep_mask;

  //recursive definition of committable elements relative to head
  //an element is committable if its rob_idx is committable and all prior elements until head are committable
  wire is_ldq1_committable_head_0;
  assign is_ldq1_committable_head_0 = isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[soc1.lsu.ldq_head]);
  wire is_ldq1_committable_head_1;
  assign is_ldq1_committable_head_1 = is_ldq1_committable_head_0 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +1) % 16]);
  wire is_ldq1_committable_head_2;
  assign is_ldq1_committable_head_2 = is_ldq1_committable_head_1 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +2) % 16]);
  wire is_ldq1_committable_head_3;
  assign is_ldq1_committable_head_3 = is_ldq1_committable_head_2 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +3) % 16]);
  wire is_ldq1_committable_head_4;
  assign is_ldq1_committable_head_4 = is_ldq1_committable_head_3 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +4) % 16]);
  wire is_ldq1_committable_head_5;
  assign is_ldq1_committable_head_5 = is_ldq1_committable_head_4 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +5) % 16]);
  wire is_ldq1_committable_head_6;
  assign is_ldq1_committable_head_6 = is_ldq1_committable_head_5 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +6) % 16]);
  wire is_ldq1_committable_head_7;
  assign is_ldq1_committable_head_7 = is_ldq1_committable_head_6 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +7) % 16]);
  wire is_ldq1_committable_head_8;
  assign is_ldq1_committable_head_8 = is_ldq1_committable_head_7 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +8) % 16]);
  wire is_ldq1_committable_head_9;
  assign is_ldq1_committable_head_9 = is_ldq1_committable_head_8 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +9) % 16]);
  wire is_ldq1_committable_head_10;
  assign is_ldq1_committable_head_10 = is_ldq1_committable_head_9 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +10) % 16]);
  wire is_ldq1_committable_head_11;
  assign is_ldq1_committable_head_11 = is_ldq1_committable_head_10 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +11) % 16]);
  wire is_ldq1_committable_head_12;
  assign is_ldq1_committable_head_12 = is_ldq1_committable_head_11 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +12) % 16]);
  wire is_ldq1_committable_head_13;
  assign is_ldq1_committable_head_13 = is_ldq1_committable_head_12 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +13) % 16]);
  wire is_ldq1_committable_head_14;
  assign is_ldq1_committable_head_14 = is_ldq1_committable_head_13 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +14) % 16]);
  wire is_ldq1_committable_head_15;
  assign is_ldq1_committable_head_15 = is_ldq1_committable_head_14 && isRobIdCommitable(soc1.core.rob.rob_head, root_id, ldq_rob_idx_1[(soc1.lsu.ldq_head +15) % 16]);

  //recursive definition of committable elements relative to head
  //an element is committable if its rob_idx is committable and all prior elements until head are committable
  wire is_ldq2_committable_head_0;
  assign is_ldq2_committable_head_0 = isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[soc2.lsu.ldq_head]);
  wire is_ldq2_committable_head_1;
  assign is_ldq2_committable_head_1 = is_ldq2_committable_head_0 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +1) % 16]);
  wire is_ldq2_committable_head_2;
  assign is_ldq2_committable_head_2 = is_ldq2_committable_head_1 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +2) % 16]);
  wire is_ldq2_committable_head_3;
  assign is_ldq2_committable_head_3 = is_ldq2_committable_head_2 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +3) % 16]);
  wire is_ldq2_committable_head_4;
  assign is_ldq2_committable_head_4 = is_ldq2_committable_head_3 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +4) % 16]);
  wire is_ldq2_committable_head_5;
  assign is_ldq2_committable_head_5 = is_ldq2_committable_head_4 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +5) % 16]);
  wire is_ldq2_committable_head_6;
  assign is_ldq2_committable_head_6 = is_ldq2_committable_head_5 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +6) % 16]);
  wire is_ldq2_committable_head_7;
  assign is_ldq2_committable_head_7 = is_ldq2_committable_head_6 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +7) % 16]);
  wire is_ldq2_committable_head_8;
  assign is_ldq2_committable_head_8 = is_ldq2_committable_head_7 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +8) % 16]);
  wire is_ldq2_committable_head_9;
  assign is_ldq2_committable_head_9 = is_ldq2_committable_head_8 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +9) % 16]);
  wire is_ldq2_committable_head_10;
  assign is_ldq2_committable_head_10 = is_ldq2_committable_head_9 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +10) % 16]);
  wire is_ldq2_committable_head_11;
  assign is_ldq2_committable_head_11 = is_ldq2_committable_head_10 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +11) % 16]);
  wire is_ldq2_committable_head_12;
  assign is_ldq2_committable_head_12 = is_ldq2_committable_head_11 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +12) % 16]);
  wire is_ldq2_committable_head_13;
  assign is_ldq2_committable_head_13 = is_ldq2_committable_head_12 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +13) % 16]);
  wire is_ldq2_committable_head_14;
  assign is_ldq2_committable_head_14 = is_ldq2_committable_head_13 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +14) % 16]);
  wire is_ldq2_committable_head_15;
  assign is_ldq2_committable_head_15 = is_ldq2_committable_head_14 && isRobIdCommitable(soc2.core.rob.rob_head, root_id, ldq_rob_idx_2[(soc2.lsu.ldq_head +15) % 16]);

  //function that maps the rob_idx to the "head-relative" entry
  function automatic is_ldq1_committable;
    //4-bit ID of the load queue entry
    input [3:0] idx;
    begin
      //mapping: (position of entry relative to head) -> (actual index of entry)
      case(idx)
        soc1.lsu.ldq_head         : is_ldq1_committable = is_ldq1_committable_head_0;
        (soc1.lsu.ldq_head+1)%16  : is_ldq1_committable = is_ldq1_committable_head_1;
        (soc1.lsu.ldq_head+2)%16  : is_ldq1_committable = is_ldq1_committable_head_2;
        (soc1.lsu.ldq_head+3)%16  : is_ldq1_committable = is_ldq1_committable_head_3;
        (soc1.lsu.ldq_head+4)%16  : is_ldq1_committable = is_ldq1_committable_head_4;
        (soc1.lsu.ldq_head+5)%16  : is_ldq1_committable = is_ldq1_committable_head_5;
        (soc1.lsu.ldq_head+6)%16  : is_ldq1_committable = is_ldq1_committable_head_6;
        (soc1.lsu.ldq_head+7)%16  : is_ldq1_committable = is_ldq1_committable_head_7;
        (soc1.lsu.ldq_head+8)%16  : is_ldq1_committable = is_ldq1_committable_head_8;
        (soc1.lsu.ldq_head+9)%16  : is_ldq1_committable = is_ldq1_committable_head_9;
        (soc1.lsu.ldq_head+10)%16 : is_ldq1_committable = is_ldq1_committable_head_10;
        (soc1.lsu.ldq_head+11)%16 : is_ldq1_committable = is_ldq1_committable_head_11;
        (soc1.lsu.ldq_head+12)%16 : is_ldq1_committable = is_ldq1_committable_head_12;
        (soc1.lsu.ldq_head+13)%16 : is_ldq1_committable = is_ldq1_committable_head_13;
        (soc1.lsu.ldq_head+14)%16 : is_ldq1_committable = is_ldq1_committable_head_14;
        (soc1.lsu.ldq_head+15)%16 : is_ldq1_committable = is_ldq1_committable_head_15;
        default                   : is_ldq1_committable = 1'b0;
      endcase
    end
  endfunction

  //function that maps the rob_idx to the "head-relative" entry
  function automatic is_ldq2_committable;
    //4-bit ID of the load queue entry
    input [3:0] idx;
    begin
      //mapping: (position of entry relative to head) -> (actual index of entry)
      case(idx)
        soc2.lsu.ldq_head         : is_ldq2_committable = is_ldq2_committable_head_0;
        (soc2.lsu.ldq_head+1)%16  : is_ldq2_committable = is_ldq2_committable_head_1;
        (soc2.lsu.ldq_head+2)%16  : is_ldq2_committable = is_ldq2_committable_head_2;
        (soc2.lsu.ldq_head+3)%16  : is_ldq2_committable = is_ldq2_committable_head_3;
        (soc2.lsu.ldq_head+4)%16  : is_ldq2_committable = is_ldq2_committable_head_4;
        (soc2.lsu.ldq_head+5)%16  : is_ldq2_committable = is_ldq2_committable_head_5;
        (soc2.lsu.ldq_head+6)%16  : is_ldq2_committable = is_ldq2_committable_head_6;
        (soc2.lsu.ldq_head+7)%16  : is_ldq2_committable = is_ldq2_committable_head_7;
        (soc2.lsu.ldq_head+8)%16  : is_ldq2_committable = is_ldq2_committable_head_8;
        (soc2.lsu.ldq_head+9)%16  : is_ldq2_committable = is_ldq2_committable_head_9;
        (soc2.lsu.ldq_head+10)%16 : is_ldq2_committable = is_ldq2_committable_head_10;
        (soc2.lsu.ldq_head+11)%16 : is_ldq2_committable = is_ldq2_committable_head_11;
        (soc2.lsu.ldq_head+12)%16 : is_ldq2_committable = is_ldq2_committable_head_12;
        (soc2.lsu.ldq_head+13)%16 : is_ldq2_committable = is_ldq2_committable_head_13;
        (soc2.lsu.ldq_head+14)%16 : is_ldq2_committable = is_ldq2_committable_head_14;
        (soc2.lsu.ldq_head+15)%16 : is_ldq2_committable = is_ldq2_committable_head_15;
        default                   : is_ldq2_committable = 1'b0;
      endcase
    end
  endfunction

	//check for all ldq entries:
	//if the entry is committable, its st_dep_mask must not overlap with the set of all uncommittable st_dep_masks
	wire st_dep_mask_consistency;
	assign st_dep_mask_consistency =
	(is_ldq1_committable(4'b0000) ? ((soc1.lsu.ldq_0_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b0001) ? ((soc1.lsu.ldq_1_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b0010) ? ((soc1.lsu.ldq_2_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b0011) ? ((soc1.lsu.ldq_3_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b0100) ? ((soc1.lsu.ldq_4_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b0101) ? ((soc1.lsu.ldq_5_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b0110) ? ((soc1.lsu.ldq_6_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b0111) ? ((soc1.lsu.ldq_7_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b1000) ? ((soc1.lsu.ldq_8_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b1001) ? ((soc1.lsu.ldq_9_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b1010) ? ((soc1.lsu.ldq_10_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b1011) ? ((soc1.lsu.ldq_11_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b1100) ? ((soc1.lsu.ldq_12_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b1101) ? ((soc1.lsu.ldq_13_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b1110) ? ((soc1.lsu.ldq_14_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq1_committable(4'b1111) ? ((soc1.lsu.ldq_15_bits_st_dep_mask & uncom1_st_dep_mask) == 16'b0) : 1'b1)  &&

	(is_ldq2_committable(4'b0000) ? ((soc2.lsu.ldq_0_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b0001) ? ((soc2.lsu.ldq_1_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b0010) ? ((soc2.lsu.ldq_2_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b0011) ? ((soc2.lsu.ldq_3_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b0100) ? ((soc2.lsu.ldq_4_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b0101) ? ((soc2.lsu.ldq_5_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b0110) ? ((soc2.lsu.ldq_6_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b0111) ? ((soc2.lsu.ldq_7_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b1000) ? ((soc2.lsu.ldq_8_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b1001) ? ((soc2.lsu.ldq_9_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b1010) ? ((soc2.lsu.ldq_10_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b1011) ? ((soc2.lsu.ldq_11_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b1100) ? ((soc2.lsu.ldq_12_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b1101) ? ((soc2.lsu.ldq_13_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b1110) ? ((soc2.lsu.ldq_14_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1)  &&
	(is_ldq2_committable(4'b1111) ? ((soc2.lsu.ldq_15_bits_st_dep_mask & uncom2_st_dep_mask) == 16'b0) : 1'b1);

  //function that returns the first uncommittable entry relative to head
  function automatic getFirstUncomLDQ1;
    begin
      case(1'b0)
        is_ldq1_committable_head_0  : getFirstUncomLDQ1 = soc1.lsu.ldq_head;
        is_ldq1_committable_head_1  : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+1)%16;
        is_ldq1_committable_head_2  : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+2)%16;
        is_ldq1_committable_head_3  : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+3)%16;
        is_ldq1_committable_head_4  : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+4)%16;
        is_ldq1_committable_head_5  : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+5)%16;
        is_ldq1_committable_head_6  : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+6)%16;
        is_ldq1_committable_head_7  : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+7)%16;
        is_ldq1_committable_head_8  : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+8)%16;
        is_ldq1_committable_head_9  : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+9)%16;
        is_ldq1_committable_head_10 : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+10)%16;
        is_ldq1_committable_head_11 : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+11)%16;
        is_ldq1_committable_head_12 : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+12)%16;
        is_ldq1_committable_head_13 : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+13)%16;
        is_ldq1_committable_head_14 : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+14)%16;
        is_ldq1_committable_head_15 : getFirstUncomLDQ1 = (soc1.lsu.ldq_head+15)%16;
        default                     : getFirstUncomLDQ1 = 4'h0;
      endcase
    end
  endfunction

  //function that returns the first uncommittable entry relative to head
  function automatic getFirstUncomLDQ2;
    begin
      case(1'b0)
        is_ldq2_committable_head_0  : getFirstUncomLDQ2 = soc2.lsu.ldq_head;
        is_ldq2_committable_head_1  : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+1)%16;
        is_ldq2_committable_head_2  : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+2)%16;
        is_ldq2_committable_head_3  : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+3)%16;
        is_ldq2_committable_head_4  : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+4)%16;
        is_ldq2_committable_head_5  : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+5)%16;
        is_ldq2_committable_head_6  : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+6)%16;
        is_ldq2_committable_head_7  : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+7)%16;
        is_ldq2_committable_head_8  : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+8)%16;
        is_ldq2_committable_head_9  : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+9)%16;
        is_ldq2_committable_head_10 : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+10)%16;
        is_ldq2_committable_head_11 : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+11)%16;
        is_ldq2_committable_head_12 : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+12)%16;
        is_ldq2_committable_head_13 : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+13)%16;
        is_ldq2_committable_head_14 : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+14)%16;
        is_ldq2_committable_head_15 : getFirstUncomLDQ2 = (soc2.lsu.ldq_head+15)%16;
        default                     : getFirstUncomLDQ2 = 4'h0;
      endcase
    end
  endfunction

  //function that returns the first uncommittable entry relative to head
  function automatic getFirstUncomSTQ1;
    begin
      case(1'b0)
        is_stq1_committable_head_0  : getFirstUncomSTQ1 = soc1.lsu.stq_head;
        is_stq1_committable_head_1  : getFirstUncomSTQ1 = (soc1.lsu.stq_head+1)%16;
        is_stq1_committable_head_2  : getFirstUncomSTQ1 = (soc1.lsu.stq_head+2)%16;
        is_stq1_committable_head_3  : getFirstUncomSTQ1 = (soc1.lsu.stq_head+3)%16;
        is_stq1_committable_head_4  : getFirstUncomSTQ1 = (soc1.lsu.stq_head+4)%16;
        is_stq1_committable_head_5  : getFirstUncomSTQ1 = (soc1.lsu.stq_head+5)%16;
        is_stq1_committable_head_6  : getFirstUncomSTQ1 = (soc1.lsu.stq_head+6)%16;
        is_stq1_committable_head_7  : getFirstUncomSTQ1 = (soc1.lsu.stq_head+7)%16;
        is_stq1_committable_head_8  : getFirstUncomSTQ1 = (soc1.lsu.stq_head+8)%16;
        is_stq1_committable_head_9  : getFirstUncomSTQ1 = (soc1.lsu.stq_head+9)%16;
        is_stq1_committable_head_10 : getFirstUncomSTQ1 = (soc1.lsu.stq_head+10)%16;
        is_stq1_committable_head_11 : getFirstUncomSTQ1 = (soc1.lsu.stq_head+11)%16;
        is_stq1_committable_head_12 : getFirstUncomSTQ1 = (soc1.lsu.stq_head+12)%16;
        is_stq1_committable_head_13 : getFirstUncomSTQ1 = (soc1.lsu.stq_head+13)%16;
        is_stq1_committable_head_14 : getFirstUncomSTQ1 = (soc1.lsu.stq_head+14)%16;
        is_stq1_committable_head_15 : getFirstUncomSTQ1 = (soc1.lsu.stq_head+15)%16;
        default                     : getFirstUncomSTQ1 = 4'h0;
      endcase
    end
  endfunction

  //function that returns the first uncommittable entry relative to head
  function automatic getFirstUncomSTQ2;
    begin
      case(1'b0)
        is_stq2_committable_head_0  : getFirstUncomSTQ2 = soc2.lsu.stq_head;
        is_stq2_committable_head_1  : getFirstUncomSTQ2 = (soc2.lsu.stq_head+1)%16;
        is_stq2_committable_head_2  : getFirstUncomSTQ2 = (soc2.lsu.stq_head+2)%16;
        is_stq2_committable_head_3  : getFirstUncomSTQ2 = (soc2.lsu.stq_head+3)%16;
        is_stq2_committable_head_4  : getFirstUncomSTQ2 = (soc2.lsu.stq_head+4)%16;
        is_stq2_committable_head_5  : getFirstUncomSTQ2 = (soc2.lsu.stq_head+5)%16;
        is_stq2_committable_head_6  : getFirstUncomSTQ2 = (soc2.lsu.stq_head+6)%16;
        is_stq2_committable_head_7  : getFirstUncomSTQ2 = (soc2.lsu.stq_head+7)%16;
        is_stq2_committable_head_8  : getFirstUncomSTQ2 = (soc2.lsu.stq_head+8)%16;
        is_stq2_committable_head_9  : getFirstUncomSTQ2 = (soc2.lsu.stq_head+9)%16;
        is_stq2_committable_head_10 : getFirstUncomSTQ2 = (soc2.lsu.stq_head+10)%16;
        is_stq2_committable_head_11 : getFirstUncomSTQ2 = (soc2.lsu.stq_head+11)%16;
        is_stq2_committable_head_12 : getFirstUncomSTQ2 = (soc2.lsu.stq_head+12)%16;
        is_stq2_committable_head_13 : getFirstUncomSTQ2 = (soc2.lsu.stq_head+13)%16;
        is_stq2_committable_head_14 : getFirstUncomSTQ2 = (soc2.lsu.stq_head+14)%16;
        is_stq2_committable_head_15 : getFirstUncomSTQ2 = (soc2.lsu.stq_head+15)%16;
        default                     : getFirstUncomSTQ2 = 4'h0;
      endcase
    end
  endfunction

  wire [3:0] ldq1_first_uncom_idx;
  assign ldq1_first_uncom_idx = getFirstUncomLDQ1();

  wire [3:0] ldq2_first_uncom_idx;
  assign ldq2_first_uncom_idx = getFirstUncomLDQ2();

  wire [3:0] stq1_first_uncom_idx;
  assign stq1_first_uncom_idx = getFirstUncomSTQ1();

  wire [3:0] stq2_first_uncom_idx;
  assign stq2_first_uncom_idx = getFirstUncomSTQ2();

  //function that returns if id1 is older than id2 with resprect to the given head of the FIFO
  function automatic isOlder(input [3:0] id1, id2, head);
    begin
      isOlder = ((id1 < id2) ^ (id1 < head) ^ (id2 < head));
    end
  endfunction

  //check for all entries:
  //if the entry is older than the first uncommittable entry: it must have a committable rob_idx
  //else: it must have an uncommittable rob_idx
  wire ldq1_consistent_rob_idx;
  assign ldq1_consistent_rob_idx = (
    (isOlder(4'h0, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_0_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_0_bits_uop_rob_idx)) &&
    (isOlder(4'h1, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_1_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_1_bits_uop_rob_idx)) &&
    (isOlder(4'h2, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_2_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_2_bits_uop_rob_idx)) &&
    (isOlder(4'h3, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_3_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_3_bits_uop_rob_idx)) &&
    (isOlder(4'h4, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_4_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_4_bits_uop_rob_idx)) &&
    (isOlder(4'h5, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_5_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_5_bits_uop_rob_idx)) &&
    (isOlder(4'h6, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_6_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_6_bits_uop_rob_idx)) &&
    (isOlder(4'h7, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_7_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_7_bits_uop_rob_idx)) &&
    (isOlder(4'h8, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_8_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_8_bits_uop_rob_idx)) &&
    (isOlder(4'h9, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_9_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_9_bits_uop_rob_idx)) &&
    (isOlder(4'ha, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_10_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_10_bits_uop_rob_idx)) &&
    (isOlder(4'hb, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_11_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_11_bits_uop_rob_idx)) &&
    (isOlder(4'hc, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_12_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_12_bits_uop_rob_idx)) &&
    (isOlder(4'hd, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_13_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_13_bits_uop_rob_idx)) &&
    (isOlder(4'he, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_14_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_14_bits_uop_rob_idx)) &&
    (isOlder(4'hf, ldq1_first_uncom_idx, soc1.lsu.ldq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_15_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.ldq_15_bits_uop_rob_idx))
    );


  //check for all entries:
  //if the entry is older than the first uncommittable entry: it must have a committable rob_idx
  //else: it must have an uncommittable rob_idx
  wire ldq2_consistent_rob_idx;
  assign ldq2_consistent_rob_idx = (
    (isOlder(4'h0, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_0_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_0_bits_uop_rob_idx)) &&
    (isOlder(4'h1, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_1_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_1_bits_uop_rob_idx)) &&
    (isOlder(4'h2, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_2_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_2_bits_uop_rob_idx)) &&
    (isOlder(4'h3, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_3_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_3_bits_uop_rob_idx)) &&
    (isOlder(4'h4, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_4_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_4_bits_uop_rob_idx)) &&
    (isOlder(4'h5, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_5_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_5_bits_uop_rob_idx)) &&
    (isOlder(4'h6, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_6_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_6_bits_uop_rob_idx)) &&
    (isOlder(4'h7, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_7_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_7_bits_uop_rob_idx)) &&
    (isOlder(4'h8, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_8_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_8_bits_uop_rob_idx)) &&
    (isOlder(4'h9, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_9_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_9_bits_uop_rob_idx)) &&
    (isOlder(4'ha, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_10_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_10_bits_uop_rob_idx)) &&
    (isOlder(4'hb, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_11_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_11_bits_uop_rob_idx)) &&
    (isOlder(4'hc, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_12_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_12_bits_uop_rob_idx)) &&
    (isOlder(4'hd, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_13_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_13_bits_uop_rob_idx)) &&
    (isOlder(4'he, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_14_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_14_bits_uop_rob_idx)) &&
    (isOlder(4'hf, ldq2_first_uncom_idx, soc2.lsu.ldq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_15_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.ldq_15_bits_uop_rob_idx))
    );

  //check for all entries:
  //if the entry is older than the first uncommittable entry: it must have a committable rob_idx
  //else: it must have an uncommittable rob_idx
  wire stq1_consistent_rob_idx;
  assign stq1_consistent_rob_idx = (
    (isOlder(4'h0, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_0_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_0_bits_uop_rob_idx)) &&
    (isOlder(4'h1, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_1_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_1_bits_uop_rob_idx)) &&
    (isOlder(4'h2, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_2_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_2_bits_uop_rob_idx)) &&
    (isOlder(4'h3, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_3_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_3_bits_uop_rob_idx)) &&
    (isOlder(4'h4, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_4_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_4_bits_uop_rob_idx)) &&
    (isOlder(4'h5, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_5_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_5_bits_uop_rob_idx)) &&
    (isOlder(4'h6, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_6_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_6_bits_uop_rob_idx)) &&
    (isOlder(4'h7, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_7_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_7_bits_uop_rob_idx)) &&
    (isOlder(4'h8, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_8_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_8_bits_uop_rob_idx)) &&
    (isOlder(4'h9, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_9_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_9_bits_uop_rob_idx)) &&
    (isOlder(4'ha, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_10_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_10_bits_uop_rob_idx)) &&
    (isOlder(4'hb, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_11_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_11_bits_uop_rob_idx)) &&
    (isOlder(4'hc, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_12_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_12_bits_uop_rob_idx)) &&
    (isOlder(4'hd, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_13_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_13_bits_uop_rob_idx)) &&
    (isOlder(4'he, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_14_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_14_bits_uop_rob_idx)) &&
    (isOlder(4'hf, stq1_first_uncom_idx, soc1.lsu.stq_head) ?
    isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_15_bits_uop_rob_idx) :
    !isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.lsu.stq_15_bits_uop_rob_idx))
    );

  //check for all entries:
  //if the entry is older than the first uncommittable entry: it must have a committable rob_idx
  //else: it must have an uncommittable rob_idx
  wire stq2_consistent_rob_idx;
  assign stq2_consistent_rob_idx = (
    (isOlder(4'h0, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_0_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_0_bits_uop_rob_idx)) &&
    (isOlder(4'h1, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_1_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_1_bits_uop_rob_idx)) &&
    (isOlder(4'h2, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_2_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_2_bits_uop_rob_idx)) &&
    (isOlder(4'h3, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_3_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_3_bits_uop_rob_idx)) &&
    (isOlder(4'h4, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_4_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_4_bits_uop_rob_idx)) &&
    (isOlder(4'h5, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_5_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_5_bits_uop_rob_idx)) &&
    (isOlder(4'h6, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_6_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_6_bits_uop_rob_idx)) &&
    (isOlder(4'h7, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_7_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_7_bits_uop_rob_idx)) &&
    (isOlder(4'h8, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_8_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_8_bits_uop_rob_idx)) &&
    (isOlder(4'h9, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_9_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_9_bits_uop_rob_idx)) &&
    (isOlder(4'ha, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_10_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_10_bits_uop_rob_idx)) &&
    (isOlder(4'hb, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_11_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_11_bits_uop_rob_idx)) &&
    (isOlder(4'hc, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_12_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_12_bits_uop_rob_idx)) &&
    (isOlder(4'hd, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_13_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_13_bits_uop_rob_idx)) &&
    (isOlder(4'he, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_14_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_14_bits_uop_rob_idx)) &&
    (isOlder(4'hf, stq2_first_uncom_idx, soc2.lsu.stq_head) ?
    isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_15_bits_uop_rob_idx) :
    !isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.lsu.stq_15_bits_uop_rob_idx))
    );

  //AND the constraints for all queues
  wire consistent_lsu_rob_idx;
  assign consistent_lsu_rob_idx = ldq1_consistent_rob_idx & ldq2_consistent_rob_idx & stq1_consistent_rob_idx & stq2_consistent_rob_idx;

      wire com_mispred_kills_root;
      assign com_mispred_kills_root =
        (mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) ?
        ((soc1.core.brinfos_0_mispredict == 1'b1) && (soc1.core.brinfos_0_valid == 1'b1) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.brinfos_0_uop_rob_idx) == 1'b1) ?
            (soc1.core.b1_mispredict_mask & root_br_mask) == root_br_mask  : 1'b1) &&
        ((soc1.core.brinfos_1_mispredict == 1'b1) && (soc1.core.brinfos_1_valid == 1'b1) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.brinfos_1_uop_rob_idx) == 1'b1) ?
            (soc1.core.b1_mispredict_mask & root_br_mask) == root_br_mask  : 1'b1) &&
        ((soc2.core.brinfos_0_mispredict == 1'b1) && (soc2.core.brinfos_0_valid == 1'b1) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.brinfos_0_uop_rob_idx) == 1'b1) ?
            (soc2.core.b1_mispredict_mask & root_br_mask) == root_br_mask  : 1'b1) &&
        ((soc2.core.brinfos_1_mispredict == 1'b1) && (soc2.core.brinfos_1_valid == 1'b1) && (isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.brinfos_1_uop_rob_idx) == 1'b1) ?
            (soc2.core.b1_mispredict_mask & root_br_mask) == root_br_mask  : 1'b1)
        :
        1'b1
      ;

	//wire enqueue_uncom_br_tags;
	//assign enqueue_uncom_br_tags =
	//(
	//  ((soc1.core.rob.io_enq_valids_0 == 1'b1) && ((isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.rob.io_enq_uops_0_rob_idx) == 1'b0) /*|| soc1.core.rob.io_enq_uops_0_rob_idx[5:1] == soc1.core.rob.rob_head*/) ?
	//  isSpawnTagGreater(soc1.core.rob.io_enq_uops_0_br_tag, commitable_masks_1) : 1'b1) &&
	//  ((soc1.core.rob.io_enq_valids_1 == 1'b1) && ((isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.rob.io_enq_uops_1_rob_idx) == 1'b0) /*|| soc1.core.rob.io_enq_uops_1_rob_idx[5:1] == soc1.core.rob.rob_head*/) ?
	//  isSpawnTagGreater(soc1.core.rob.io_enq_uops_1_br_tag, commitable_masks_1) : 1'b1) &&
	//  ((soc2.core.rob.io_enq_valids_0 == 1'b1) && ((isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.rob.io_enq_uops_0_rob_idx) == 1'b0) /*|| soc2.core.rob.io_enq_uops_0_rob_idx[5:1] == soc2.core.rob.rob_head*/) ?
	//  isSpawnTagGreater(soc2.core.rob.io_enq_uops_0_br_tag, commitable_masks_2) : 1'b1) &&
	//  ((soc2.core.rob.io_enq_valids_1 == 1'b1) && ((isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.rob.io_enq_uops_1_rob_idx) == 1'b0) /*|| soc2.core.rob.io_enq_uops_1_rob_idx[5:1] == soc2.core.rob.rob_head*/) ?
	//  isSpawnTagGreater(soc2.core.rob.io_enq_uops_1_br_tag, commitable_masks_2) : 1'b1)
	//);

	//check for all ROB entries:
	//if entry is older than tail and younger than root_id
	//its branch mask must contain root_br_mask and it is valid
	//or the entry is invalid
	wire consistent_uncommittable_masks;
	assign consistent_uncommittable_masks =
	  (!mispred_happened_1 && !mispred_happened_2 && !root_id_killed && !root_id_already_killed)
	  ? 
	  (ROBisOlder(6'h0,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h0] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h0] == 1'b1)) || (rob_valids_1[6'h0] == 1'b0) : (((rob_branch_masks_1[6'h0] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h0] == 1'b1)) || (rob_valids_1[6'h0] == 1'b0)) &&
	  (ROBisOlder(6'h1,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h1] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h1] == 1'b1)) || (rob_valids_1[6'h1] == 1'b0) : (((rob_branch_masks_1[6'h1] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h1] == 1'b1)) || (rob_valids_1[6'h1] == 1'b0)) &&
	  (ROBisOlder(6'h2,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h2] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h2] == 1'b1)) || (rob_valids_1[6'h2] == 1'b0) : (((rob_branch_masks_1[6'h2] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h2] == 1'b1)) || (rob_valids_1[6'h2] == 1'b0)) &&
	  (ROBisOlder(6'h3,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h3] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h3] == 1'b1)) || (rob_valids_1[6'h3] == 1'b0) : (((rob_branch_masks_1[6'h3] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h3] == 1'b1)) || (rob_valids_1[6'h3] == 1'b0)) &&
	  (ROBisOlder(6'h4,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h4] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h4] == 1'b1)) || (rob_valids_1[6'h4] == 1'b0) : (((rob_branch_masks_1[6'h4] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h4] == 1'b1)) || (rob_valids_1[6'h4] == 1'b0)) &&
	  (ROBisOlder(6'h5,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h5] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h5] == 1'b1)) || (rob_valids_1[6'h5] == 1'b0) : (((rob_branch_masks_1[6'h5] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h5] == 1'b1)) || (rob_valids_1[6'h5] == 1'b0)) &&
	  (ROBisOlder(6'h6,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h6] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h6] == 1'b1)) || (rob_valids_1[6'h6] == 1'b0) : (((rob_branch_masks_1[6'h6] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h6] == 1'b1)) || (rob_valids_1[6'h6] == 1'b0)) &&
	  (ROBisOlder(6'h7,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h7] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h7] == 1'b1)) || (rob_valids_1[6'h7] == 1'b0) : (((rob_branch_masks_1[6'h7] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h7] == 1'b1)) || (rob_valids_1[6'h7] == 1'b0)) &&
	  (ROBisOlder(6'h8,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h8] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h8] == 1'b1)) || (rob_valids_1[6'h8] == 1'b0) : (((rob_branch_masks_1[6'h8] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h8] == 1'b1)) || (rob_valids_1[6'h8] == 1'b0)) &&
	  (ROBisOlder(6'h9,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h9] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h9] == 1'b1)) || (rob_valids_1[6'h9] == 1'b0) : (((rob_branch_masks_1[6'h9] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h9] == 1'b1)) || (rob_valids_1[6'h9] == 1'b0)) &&
	  (ROBisOlder(6'ha,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'ha] & root_br_mask) == root_br_mask) && (rob_valids_1[6'ha] == 1'b1)) || (rob_valids_1[6'ha] == 1'b0) : (((rob_branch_masks_1[6'ha] & root_br_mask) != root_br_mask) && (rob_valids_1[6'ha] == 1'b1)) || (rob_valids_1[6'ha] == 1'b0)) &&
	  (ROBisOlder(6'hb,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'hb] & root_br_mask) == root_br_mask) && (rob_valids_1[6'hb] == 1'b1)) || (rob_valids_1[6'hb] == 1'b0) : (((rob_branch_masks_1[6'hb] & root_br_mask) != root_br_mask) && (rob_valids_1[6'hb] == 1'b1)) || (rob_valids_1[6'hb] == 1'b0)) &&
	  (ROBisOlder(6'hc,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'hc] & root_br_mask) == root_br_mask) && (rob_valids_1[6'hc] == 1'b1)) || (rob_valids_1[6'hc] == 1'b0) : (((rob_branch_masks_1[6'hc] & root_br_mask) != root_br_mask) && (rob_valids_1[6'hc] == 1'b1)) || (rob_valids_1[6'hc] == 1'b0)) &&
	  (ROBisOlder(6'hd,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'hd] & root_br_mask) == root_br_mask) && (rob_valids_1[6'hd] == 1'b1)) || (rob_valids_1[6'hd] == 1'b0) : (((rob_branch_masks_1[6'hd] & root_br_mask) != root_br_mask) && (rob_valids_1[6'hd] == 1'b1)) || (rob_valids_1[6'hd] == 1'b0)) &&
	  (ROBisOlder(6'he,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'he] & root_br_mask) == root_br_mask) && (rob_valids_1[6'he] == 1'b1)) || (rob_valids_1[6'he] == 1'b0) : (((rob_branch_masks_1[6'he] & root_br_mask) != root_br_mask) && (rob_valids_1[6'he] == 1'b1)) || (rob_valids_1[6'he] == 1'b0)) &&
	  (ROBisOlder(6'hf,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'hf] & root_br_mask) == root_br_mask) && (rob_valids_1[6'hf] == 1'b1)) || (rob_valids_1[6'hf] == 1'b0) : (((rob_branch_masks_1[6'hf] & root_br_mask) != root_br_mask) && (rob_valids_1[6'hf] == 1'b1)) || (rob_valids_1[6'hf] == 1'b0)) &&
	  (ROBisOlder(6'h10,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h10] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h10] == 1'b1)) || (rob_valids_1[6'h10] == 1'b0) : (((rob_branch_masks_1[6'h10] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h10] == 1'b1)) || (rob_valids_1[6'h10] == 1'b0)) &&
	  (ROBisOlder(6'h11,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h11] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h11] == 1'b1)) || (rob_valids_1[6'h11] == 1'b0) : (((rob_branch_masks_1[6'h11] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h11] == 1'b1)) || (rob_valids_1[6'h11] == 1'b0)) &&
	  (ROBisOlder(6'h12,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h12] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h12] == 1'b1)) || (rob_valids_1[6'h12] == 1'b0) : (((rob_branch_masks_1[6'h12] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h12] == 1'b1)) || (rob_valids_1[6'h12] == 1'b0)) &&
	  (ROBisOlder(6'h13,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h13] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h13] == 1'b1)) || (rob_valids_1[6'h13] == 1'b0) : (((rob_branch_masks_1[6'h13] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h13] == 1'b1)) || (rob_valids_1[6'h13] == 1'b0)) &&
	  (ROBisOlder(6'h14,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h14] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h14] == 1'b1)) || (rob_valids_1[6'h14] == 1'b0) : (((rob_branch_masks_1[6'h14] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h14] == 1'b1)) || (rob_valids_1[6'h14] == 1'b0)) &&
	  (ROBisOlder(6'h15,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h15] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h15] == 1'b1)) || (rob_valids_1[6'h15] == 1'b0) : (((rob_branch_masks_1[6'h15] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h15] == 1'b1)) || (rob_valids_1[6'h15] == 1'b0)) &&
	  (ROBisOlder(6'h16,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h16] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h16] == 1'b1)) || (rob_valids_1[6'h16] == 1'b0) : (((rob_branch_masks_1[6'h16] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h16] == 1'b1)) || (rob_valids_1[6'h16] == 1'b0)) &&
	  (ROBisOlder(6'h17,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h17] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h17] == 1'b1)) || (rob_valids_1[6'h17] == 1'b0) : (((rob_branch_masks_1[6'h17] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h17] == 1'b1)) || (rob_valids_1[6'h17] == 1'b0)) &&
	  (ROBisOlder(6'h18,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h18] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h18] == 1'b1)) || (rob_valids_1[6'h18] == 1'b0) : (((rob_branch_masks_1[6'h18] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h18] == 1'b1)) || (rob_valids_1[6'h18] == 1'b0)) &&
	  (ROBisOlder(6'h19,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h19] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h19] == 1'b1)) || (rob_valids_1[6'h19] == 1'b0) : (((rob_branch_masks_1[6'h19] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h19] == 1'b1)) || (rob_valids_1[6'h19] == 1'b0)) &&
	  (ROBisOlder(6'h1a,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h1a] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h1a] == 1'b1)) || (rob_valids_1[6'h1a] == 1'b0) : (((rob_branch_masks_1[6'h1a] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h1a] == 1'b1)) || (rob_valids_1[6'h1a] == 1'b0)) &&
	  (ROBisOlder(6'h1b,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h1b] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h1b] == 1'b1)) || (rob_valids_1[6'h1b] == 1'b0) : (((rob_branch_masks_1[6'h1b] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h1b] == 1'b1)) || (rob_valids_1[6'h1b] == 1'b0)) &&
	  (ROBisOlder(6'h1c,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h1c] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h1c] == 1'b1)) || (rob_valids_1[6'h1c] == 1'b0) : (((rob_branch_masks_1[6'h1c] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h1c] == 1'b1)) || (rob_valids_1[6'h1c] == 1'b0)) &&
	  (ROBisOlder(6'h1d,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h1d] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h1d] == 1'b1)) || (rob_valids_1[6'h1d] == 1'b0) : (((rob_branch_masks_1[6'h1d] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h1d] == 1'b1)) || (rob_valids_1[6'h1d] == 1'b0)) &&
	  (ROBisOlder(6'h1e,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h1e] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h1e] == 1'b1)) || (rob_valids_1[6'h1e] == 1'b0) : (((rob_branch_masks_1[6'h1e] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h1e] == 1'b1)) || (rob_valids_1[6'h1e] == 1'b0)) &&
	  (ROBisOlder(6'h1f,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h1f] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h1f] == 1'b1)) || (rob_valids_1[6'h1f] == 1'b0) : (((rob_branch_masks_1[6'h1f] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h1f] == 1'b1)) || (rob_valids_1[6'h1f] == 1'b0)) &&
	  (ROBisOlder(6'h20,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h20] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h20] == 1'b1)) || (rob_valids_1[6'h20] == 1'b0) : (((rob_branch_masks_1[6'h20] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h20] == 1'b1)) || (rob_valids_1[6'h20] == 1'b0)) &&
	  (ROBisOlder(6'h21,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h21] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h21] == 1'b1)) || (rob_valids_1[6'h21] == 1'b0) : (((rob_branch_masks_1[6'h21] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h21] == 1'b1)) || (rob_valids_1[6'h21] == 1'b0)) &&
	  (ROBisOlder(6'h22,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h22] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h22] == 1'b1)) || (rob_valids_1[6'h22] == 1'b0) : (((rob_branch_masks_1[6'h22] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h22] == 1'b1)) || (rob_valids_1[6'h22] == 1'b0)) &&
	  (ROBisOlder(6'h23,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h23] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h23] == 1'b1)) || (rob_valids_1[6'h23] == 1'b0) : (((rob_branch_masks_1[6'h23] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h23] == 1'b1)) || (rob_valids_1[6'h23] == 1'b0)) &&
	  (ROBisOlder(6'h24,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h24] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h24] == 1'b1)) || (rob_valids_1[6'h24] == 1'b0) : (((rob_branch_masks_1[6'h24] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h24] == 1'b1)) || (rob_valids_1[6'h24] == 1'b0)) &&
	  (ROBisOlder(6'h25,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h25] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h25] == 1'b1)) || (rob_valids_1[6'h25] == 1'b0) : (((rob_branch_masks_1[6'h25] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h25] == 1'b1)) || (rob_valids_1[6'h25] == 1'b0)) &&
	  (ROBisOlder(6'h26,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h26] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h26] == 1'b1)) || (rob_valids_1[6'h26] == 1'b0) : (((rob_branch_masks_1[6'h26] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h26] == 1'b1)) || (rob_valids_1[6'h26] == 1'b0)) &&
	  (ROBisOlder(6'h27,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h27] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h27] == 1'b1)) || (rob_valids_1[6'h27] == 1'b0) : (((rob_branch_masks_1[6'h27] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h27] == 1'b1)) || (rob_valids_1[6'h27] == 1'b0)) &&
	  (ROBisOlder(6'h28,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h28] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h28] == 1'b1)) || (rob_valids_1[6'h28] == 1'b0) : (((rob_branch_masks_1[6'h28] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h28] == 1'b1)) || (rob_valids_1[6'h28] == 1'b0)) &&
	  (ROBisOlder(6'h29,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h29] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h29] == 1'b1)) || (rob_valids_1[6'h29] == 1'b0) : (((rob_branch_masks_1[6'h29] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h29] == 1'b1)) || (rob_valids_1[6'h29] == 1'b0)) &&
	  (ROBisOlder(6'h2a,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h2a] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h2a] == 1'b1)) || (rob_valids_1[6'h2a] == 1'b0) : (((rob_branch_masks_1[6'h2a] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h2a] == 1'b1)) || (rob_valids_1[6'h2a] == 1'b0)) &&
	  (ROBisOlder(6'h2b,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h2b] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h2b] == 1'b1)) || (rob_valids_1[6'h2b] == 1'b0) : (((rob_branch_masks_1[6'h2b] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h2b] == 1'b1)) || (rob_valids_1[6'h2b] == 1'b0)) &&
	  (ROBisOlder(6'h2c,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h2c] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h2c] == 1'b1)) || (rob_valids_1[6'h2c] == 1'b0) : (((rob_branch_masks_1[6'h2c] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h2c] == 1'b1)) || (rob_valids_1[6'h2c] == 1'b0)) &&
	  (ROBisOlder(6'h2d,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h2d] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h2d] == 1'b1)) || (rob_valids_1[6'h2d] == 1'b0) : (((rob_branch_masks_1[6'h2d] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h2d] == 1'b1)) || (rob_valids_1[6'h2d] == 1'b0)) &&
	  (ROBisOlder(6'h2e,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h2e] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h2e] == 1'b1)) || (rob_valids_1[6'h2e] == 1'b0) : (((rob_branch_masks_1[6'h2e] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h2e] == 1'b1)) || (rob_valids_1[6'h2e] == 1'b0)) &&
	  (ROBisOlder(6'h2f,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h2f] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h2f] == 1'b1)) || (rob_valids_1[6'h2f] == 1'b0) : (((rob_branch_masks_1[6'h2f] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h2f] == 1'b1)) || (rob_valids_1[6'h2f] == 1'b0)) &&
	  (ROBisOlder(6'h30,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h30] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h30] == 1'b1)) || (rob_valids_1[6'h30] == 1'b0) : (((rob_branch_masks_1[6'h30] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h30] == 1'b1)) || (rob_valids_1[6'h30] == 1'b0)) &&
	  (ROBisOlder(6'h31,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h31] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h31] == 1'b1)) || (rob_valids_1[6'h31] == 1'b0) : (((rob_branch_masks_1[6'h31] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h31] == 1'b1)) || (rob_valids_1[6'h31] == 1'b0)) &&
	  (ROBisOlder(6'h32,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h32] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h32] == 1'b1)) || (rob_valids_1[6'h32] == 1'b0) : (((rob_branch_masks_1[6'h32] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h32] == 1'b1)) || (rob_valids_1[6'h32] == 1'b0)) &&
	  (ROBisOlder(6'h33,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h33] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h33] == 1'b1)) || (rob_valids_1[6'h33] == 1'b0) : (((rob_branch_masks_1[6'h33] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h33] == 1'b1)) || (rob_valids_1[6'h33] == 1'b0)) &&
	  (ROBisOlder(6'h34,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h34] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h34] == 1'b1)) || (rob_valids_1[6'h34] == 1'b0) : (((rob_branch_masks_1[6'h34] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h34] == 1'b1)) || (rob_valids_1[6'h34] == 1'b0)) &&
	  (ROBisOlder(6'h35,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h35] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h35] == 1'b1)) || (rob_valids_1[6'h35] == 1'b0) : (((rob_branch_masks_1[6'h35] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h35] == 1'b1)) || (rob_valids_1[6'h35] == 1'b0)) &&
	  (ROBisOlder(6'h36,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h36] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h36] == 1'b1)) || (rob_valids_1[6'h36] == 1'b0) : (((rob_branch_masks_1[6'h36] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h36] == 1'b1)) || (rob_valids_1[6'h36] == 1'b0)) &&
	  (ROBisOlder(6'h37,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h37] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h37] == 1'b1)) || (rob_valids_1[6'h37] == 1'b0) : (((rob_branch_masks_1[6'h37] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h37] == 1'b1)) || (rob_valids_1[6'h37] == 1'b0)) &&
	  (ROBisOlder(6'h38,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h38] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h38] == 1'b1)) || (rob_valids_1[6'h38] == 1'b0) : (((rob_branch_masks_1[6'h38] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h38] == 1'b1)) || (rob_valids_1[6'h38] == 1'b0)) &&
	  (ROBisOlder(6'h39,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h39] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h39] == 1'b1)) || (rob_valids_1[6'h39] == 1'b0) : (((rob_branch_masks_1[6'h39] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h39] == 1'b1)) || (rob_valids_1[6'h39] == 1'b0)) &&
	  (ROBisOlder(6'h3a,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h3a] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h3a] == 1'b1)) || (rob_valids_1[6'h3a] == 1'b0) : (((rob_branch_masks_1[6'h3a] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h3a] == 1'b1)) || (rob_valids_1[6'h3a] == 1'b0)) &&
	  (ROBisOlder(6'h3b,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h3b] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h3b] == 1'b1)) || (rob_valids_1[6'h3b] == 1'b0) : (((rob_branch_masks_1[6'h3b] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h3b] == 1'b1)) || (rob_valids_1[6'h3b] == 1'b0)) &&
	  (ROBisOlder(6'h3c,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h3c] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h3c] == 1'b1)) || (rob_valids_1[6'h3c] == 1'b0) : (((rob_branch_masks_1[6'h3c] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h3c] == 1'b1)) || (rob_valids_1[6'h3c] == 1'b0)) &&
	  (ROBisOlder(6'h3d,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h3d] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h3d] == 1'b1)) || (rob_valids_1[6'h3d] == 1'b0) : (((rob_branch_masks_1[6'h3d] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h3d] == 1'b1)) || (rob_valids_1[6'h3d] == 1'b0)) &&
	  (ROBisOlder(6'h3e,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h3e] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h3e] == 1'b1)) || (rob_valids_1[6'h3e] == 1'b0) : (((rob_branch_masks_1[6'h3e] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h3e] == 1'b1)) || (rob_valids_1[6'h3e] == 1'b0)) &&
	  (ROBisOlder(6'h3f,soc1.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_1[6'h3f] & root_br_mask) == root_br_mask) && (rob_valids_1[6'h3f] == 1'b1)) || (rob_valids_1[6'h3f] == 1'b0) : (((rob_branch_masks_1[6'h3f] & root_br_mask) != root_br_mask) && (rob_valids_1[6'h3f] == 1'b1)) || (rob_valids_1[6'h3f] == 1'b0)) &&

	  (ROBisOlder(6'h0,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h0] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h0] == 1'b1)) || (rob_valids_2[6'h0] == 1'b0) : (((rob_branch_masks_2[6'h0] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h0] == 1'b1)) || (rob_valids_2[6'h0] == 1'b0)) &&
	  (ROBisOlder(6'h1,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h1] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h1] == 1'b1)) || (rob_valids_2[6'h1] == 1'b0) : (((rob_branch_masks_2[6'h1] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h1] == 1'b1)) || (rob_valids_2[6'h1] == 1'b0)) &&
	  (ROBisOlder(6'h2,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h2] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h2] == 1'b1)) || (rob_valids_2[6'h2] == 1'b0) : (((rob_branch_masks_2[6'h2] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h2] == 1'b1)) || (rob_valids_2[6'h2] == 1'b0)) &&
	  (ROBisOlder(6'h3,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h3] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h3] == 1'b1)) || (rob_valids_2[6'h3] == 1'b0) : (((rob_branch_masks_2[6'h3] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h3] == 1'b1)) || (rob_valids_2[6'h3] == 1'b0)) &&
	  (ROBisOlder(6'h4,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h4] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h4] == 1'b1)) || (rob_valids_2[6'h4] == 1'b0) : (((rob_branch_masks_2[6'h4] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h4] == 1'b1)) || (rob_valids_2[6'h4] == 1'b0)) &&
	  (ROBisOlder(6'h5,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h5] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h5] == 1'b1)) || (rob_valids_2[6'h5] == 1'b0) : (((rob_branch_masks_2[6'h5] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h5] == 1'b1)) || (rob_valids_2[6'h5] == 1'b0)) &&
	  (ROBisOlder(6'h6,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h6] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h6] == 1'b1)) || (rob_valids_2[6'h6] == 1'b0) : (((rob_branch_masks_2[6'h6] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h6] == 1'b1)) || (rob_valids_2[6'h6] == 1'b0)) &&
	  (ROBisOlder(6'h7,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h7] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h7] == 1'b1)) || (rob_valids_2[6'h7] == 1'b0) : (((rob_branch_masks_2[6'h7] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h7] == 1'b1)) || (rob_valids_2[6'h7] == 1'b0)) &&
	  (ROBisOlder(6'h8,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h8] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h8] == 1'b1)) || (rob_valids_2[6'h8] == 1'b0) : (((rob_branch_masks_2[6'h8] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h8] == 1'b1)) || (rob_valids_2[6'h8] == 1'b0)) &&
	  (ROBisOlder(6'h9,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h9] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h9] == 1'b1)) || (rob_valids_2[6'h9] == 1'b0) : (((rob_branch_masks_2[6'h9] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h9] == 1'b1)) || (rob_valids_2[6'h9] == 1'b0)) &&
	  (ROBisOlder(6'ha,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'ha] & root_br_mask) == root_br_mask) && (rob_valids_2[6'ha] == 1'b1)) || (rob_valids_2[6'ha] == 1'b0) : (((rob_branch_masks_2[6'ha] & root_br_mask) != root_br_mask) && (rob_valids_2[6'ha] == 1'b1)) || (rob_valids_2[6'ha] == 1'b0)) &&
	  (ROBisOlder(6'hb,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'hb] & root_br_mask) == root_br_mask) && (rob_valids_2[6'hb] == 1'b1)) || (rob_valids_2[6'hb] == 1'b0) : (((rob_branch_masks_2[6'hb] & root_br_mask) != root_br_mask) && (rob_valids_2[6'hb] == 1'b1)) || (rob_valids_2[6'hb] == 1'b0)) &&
	  (ROBisOlder(6'hc,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'hc] & root_br_mask) == root_br_mask) && (rob_valids_2[6'hc] == 1'b1)) || (rob_valids_2[6'hc] == 1'b0) : (((rob_branch_masks_2[6'hc] & root_br_mask) != root_br_mask) && (rob_valids_2[6'hc] == 1'b1)) || (rob_valids_2[6'hc] == 1'b0)) &&
	  (ROBisOlder(6'hd,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'hd] & root_br_mask) == root_br_mask) && (rob_valids_2[6'hd] == 1'b1)) || (rob_valids_2[6'hd] == 1'b0) : (((rob_branch_masks_2[6'hd] & root_br_mask) != root_br_mask) && (rob_valids_2[6'hd] == 1'b1)) || (rob_valids_2[6'hd] == 1'b0)) &&
	  (ROBisOlder(6'he,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'he] & root_br_mask) == root_br_mask) && (rob_valids_2[6'he] == 1'b1)) || (rob_valids_2[6'he] == 1'b0) : (((rob_branch_masks_2[6'he] & root_br_mask) != root_br_mask) && (rob_valids_2[6'he] == 1'b1)) || (rob_valids_2[6'he] == 1'b0)) &&
	  (ROBisOlder(6'hf,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'hf] & root_br_mask) == root_br_mask) && (rob_valids_2[6'hf] == 1'b1)) || (rob_valids_2[6'hf] == 1'b0) : (((rob_branch_masks_2[6'hf] & root_br_mask) != root_br_mask) && (rob_valids_2[6'hf] == 1'b1)) || (rob_valids_2[6'hf] == 1'b0)) &&
	  (ROBisOlder(6'h10,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h10] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h10] == 1'b1)) || (rob_valids_2[6'h10] == 1'b0) : (((rob_branch_masks_2[6'h10] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h10] == 1'b1)) || (rob_valids_2[6'h10] == 1'b0)) &&
	  (ROBisOlder(6'h11,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h11] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h11] == 1'b1)) || (rob_valids_2[6'h11] == 1'b0) : (((rob_branch_masks_2[6'h11] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h11] == 1'b1)) || (rob_valids_2[6'h11] == 1'b0)) &&
	  (ROBisOlder(6'h12,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h12] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h12] == 1'b1)) || (rob_valids_2[6'h12] == 1'b0) : (((rob_branch_masks_2[6'h12] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h12] == 1'b1)) || (rob_valids_2[6'h12] == 1'b0)) &&
	  (ROBisOlder(6'h13,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h13] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h13] == 1'b1)) || (rob_valids_2[6'h13] == 1'b0) : (((rob_branch_masks_2[6'h13] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h13] == 1'b1)) || (rob_valids_2[6'h13] == 1'b0)) &&
	  (ROBisOlder(6'h14,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h14] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h14] == 1'b1)) || (rob_valids_2[6'h14] == 1'b0) : (((rob_branch_masks_2[6'h14] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h14] == 1'b1)) || (rob_valids_2[6'h14] == 1'b0)) &&
	  (ROBisOlder(6'h15,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h15] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h15] == 1'b1)) || (rob_valids_2[6'h15] == 1'b0) : (((rob_branch_masks_2[6'h15] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h15] == 1'b1)) || (rob_valids_2[6'h15] == 1'b0)) &&
	  (ROBisOlder(6'h16,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h16] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h16] == 1'b1)) || (rob_valids_2[6'h16] == 1'b0) : (((rob_branch_masks_2[6'h16] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h16] == 1'b1)) || (rob_valids_2[6'h16] == 1'b0)) &&
	  (ROBisOlder(6'h17,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h17] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h17] == 1'b1)) || (rob_valids_2[6'h17] == 1'b0) : (((rob_branch_masks_2[6'h17] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h17] == 1'b1)) || (rob_valids_2[6'h17] == 1'b0)) &&
	  (ROBisOlder(6'h18,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h18] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h18] == 1'b1)) || (rob_valids_2[6'h18] == 1'b0) : (((rob_branch_masks_2[6'h18] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h18] == 1'b1)) || (rob_valids_2[6'h18] == 1'b0)) &&
	  (ROBisOlder(6'h19,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h19] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h19] == 1'b1)) || (rob_valids_2[6'h19] == 1'b0) : (((rob_branch_masks_2[6'h19] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h19] == 1'b1)) || (rob_valids_2[6'h19] == 1'b0)) &&
	  (ROBisOlder(6'h1a,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h1a] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h1a] == 1'b1)) || (rob_valids_2[6'h1a] == 1'b0) : (((rob_branch_masks_2[6'h1a] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h1a] == 1'b1)) || (rob_valids_2[6'h1a] == 1'b0)) &&
	  (ROBisOlder(6'h1b,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h1b] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h1b] == 1'b1)) || (rob_valids_2[6'h1b] == 1'b0) : (((rob_branch_masks_2[6'h1b] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h1b] == 1'b1)) || (rob_valids_2[6'h1b] == 1'b0)) &&
	  (ROBisOlder(6'h1c,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h1c] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h1c] == 1'b1)) || (rob_valids_2[6'h1c] == 1'b0) : (((rob_branch_masks_2[6'h1c] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h1c] == 1'b1)) || (rob_valids_2[6'h1c] == 1'b0)) &&
	  (ROBisOlder(6'h1d,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h1d] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h1d] == 1'b1)) || (rob_valids_2[6'h1d] == 1'b0) : (((rob_branch_masks_2[6'h1d] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h1d] == 1'b1)) || (rob_valids_2[6'h1d] == 1'b0)) &&
	  (ROBisOlder(6'h1e,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h1e] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h1e] == 1'b1)) || (rob_valids_2[6'h1e] == 1'b0) : (((rob_branch_masks_2[6'h1e] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h1e] == 1'b1)) || (rob_valids_2[6'h1e] == 1'b0)) &&
	  (ROBisOlder(6'h1f,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h1f] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h1f] == 1'b1)) || (rob_valids_2[6'h1f] == 1'b0) : (((rob_branch_masks_2[6'h1f] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h1f] == 1'b1)) || (rob_valids_2[6'h1f] == 1'b0)) &&
	  (ROBisOlder(6'h20,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h20] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h20] == 1'b1)) || (rob_valids_2[6'h20] == 1'b0) : (((rob_branch_masks_2[6'h20] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h20] == 1'b1)) || (rob_valids_2[6'h20] == 1'b0)) &&
	  (ROBisOlder(6'h21,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h21] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h21] == 1'b1)) || (rob_valids_2[6'h21] == 1'b0) : (((rob_branch_masks_2[6'h21] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h21] == 1'b1)) || (rob_valids_2[6'h21] == 1'b0)) &&
	  (ROBisOlder(6'h22,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h22] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h22] == 1'b1)) || (rob_valids_2[6'h22] == 1'b0) : (((rob_branch_masks_2[6'h22] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h22] == 1'b1)) || (rob_valids_2[6'h22] == 1'b0)) &&
	  (ROBisOlder(6'h23,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h23] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h23] == 1'b1)) || (rob_valids_2[6'h23] == 1'b0) : (((rob_branch_masks_2[6'h23] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h23] == 1'b1)) || (rob_valids_2[6'h23] == 1'b0)) &&
	  (ROBisOlder(6'h24,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h24] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h24] == 1'b1)) || (rob_valids_2[6'h24] == 1'b0) : (((rob_branch_masks_2[6'h24] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h24] == 1'b1)) || (rob_valids_2[6'h24] == 1'b0)) &&
	  (ROBisOlder(6'h25,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h25] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h25] == 1'b1)) || (rob_valids_2[6'h25] == 1'b0) : (((rob_branch_masks_2[6'h25] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h25] == 1'b1)) || (rob_valids_2[6'h25] == 1'b0)) &&
	  (ROBisOlder(6'h26,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h26] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h26] == 1'b1)) || (rob_valids_2[6'h26] == 1'b0) : (((rob_branch_masks_2[6'h26] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h26] == 1'b1)) || (rob_valids_2[6'h26] == 1'b0)) &&
	  (ROBisOlder(6'h27,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h27] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h27] == 1'b1)) || (rob_valids_2[6'h27] == 1'b0) : (((rob_branch_masks_2[6'h27] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h27] == 1'b1)) || (rob_valids_2[6'h27] == 1'b0)) &&
	  (ROBisOlder(6'h28,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h28] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h28] == 1'b1)) || (rob_valids_2[6'h28] == 1'b0) : (((rob_branch_masks_2[6'h28] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h28] == 1'b1)) || (rob_valids_2[6'h28] == 1'b0)) &&
	  (ROBisOlder(6'h29,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h29] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h29] == 1'b1)) || (rob_valids_2[6'h29] == 1'b0) : (((rob_branch_masks_2[6'h29] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h29] == 1'b1)) || (rob_valids_2[6'h29] == 1'b0)) &&
	  (ROBisOlder(6'h2a,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h2a] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h2a] == 1'b1)) || (rob_valids_2[6'h2a] == 1'b0) : (((rob_branch_masks_2[6'h2a] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h2a] == 1'b1)) || (rob_valids_2[6'h2a] == 1'b0)) &&
	  (ROBisOlder(6'h2b,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h2b] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h2b] == 1'b1)) || (rob_valids_2[6'h2b] == 1'b0) : (((rob_branch_masks_2[6'h2b] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h2b] == 1'b1)) || (rob_valids_2[6'h2b] == 1'b0)) &&
	  (ROBisOlder(6'h2c,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h2c] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h2c] == 1'b1)) || (rob_valids_2[6'h2c] == 1'b0) : (((rob_branch_masks_2[6'h2c] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h2c] == 1'b1)) || (rob_valids_2[6'h2c] == 1'b0)) &&
	  (ROBisOlder(6'h2d,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h2d] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h2d] == 1'b1)) || (rob_valids_2[6'h2d] == 1'b0) : (((rob_branch_masks_2[6'h2d] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h2d] == 1'b1)) || (rob_valids_2[6'h2d] == 1'b0)) &&
	  (ROBisOlder(6'h2e,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h2e] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h2e] == 1'b1)) || (rob_valids_2[6'h2e] == 1'b0) : (((rob_branch_masks_2[6'h2e] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h2e] == 1'b1)) || (rob_valids_2[6'h2e] == 1'b0)) &&
	  (ROBisOlder(6'h2f,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h2f] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h2f] == 1'b1)) || (rob_valids_2[6'h2f] == 1'b0) : (((rob_branch_masks_2[6'h2f] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h2f] == 1'b1)) || (rob_valids_2[6'h2f] == 1'b0)) &&
	  (ROBisOlder(6'h30,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h30] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h30] == 1'b1)) || (rob_valids_2[6'h30] == 1'b0) : (((rob_branch_masks_2[6'h30] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h30] == 1'b1)) || (rob_valids_2[6'h30] == 1'b0)) &&
	  (ROBisOlder(6'h31,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h31] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h31] == 1'b1)) || (rob_valids_2[6'h31] == 1'b0) : (((rob_branch_masks_2[6'h31] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h31] == 1'b1)) || (rob_valids_2[6'h31] == 1'b0)) &&
	  (ROBisOlder(6'h32,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h32] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h32] == 1'b1)) || (rob_valids_2[6'h32] == 1'b0) : (((rob_branch_masks_2[6'h32] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h32] == 1'b1)) || (rob_valids_2[6'h32] == 1'b0)) &&
	  (ROBisOlder(6'h33,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h33] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h33] == 1'b1)) || (rob_valids_2[6'h33] == 1'b0) : (((rob_branch_masks_2[6'h33] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h33] == 1'b1)) || (rob_valids_2[6'h33] == 1'b0)) &&
	  (ROBisOlder(6'h34,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h34] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h34] == 1'b1)) || (rob_valids_2[6'h34] == 1'b0) : (((rob_branch_masks_2[6'h34] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h34] == 1'b1)) || (rob_valids_2[6'h34] == 1'b0)) &&
	  (ROBisOlder(6'h35,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h35] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h35] == 1'b1)) || (rob_valids_2[6'h35] == 1'b0) : (((rob_branch_masks_2[6'h35] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h35] == 1'b1)) || (rob_valids_2[6'h35] == 1'b0)) &&
	  (ROBisOlder(6'h36,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h36] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h36] == 1'b1)) || (rob_valids_2[6'h36] == 1'b0) : (((rob_branch_masks_2[6'h36] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h36] == 1'b1)) || (rob_valids_2[6'h36] == 1'b0)) &&
	  (ROBisOlder(6'h37,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h37] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h37] == 1'b1)) || (rob_valids_2[6'h37] == 1'b0) : (((rob_branch_masks_2[6'h37] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h37] == 1'b1)) || (rob_valids_2[6'h37] == 1'b0)) &&
	  (ROBisOlder(6'h38,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h38] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h38] == 1'b1)) || (rob_valids_2[6'h38] == 1'b0) : (((rob_branch_masks_2[6'h38] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h38] == 1'b1)) || (rob_valids_2[6'h38] == 1'b0)) &&
	  (ROBisOlder(6'h39,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h39] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h39] == 1'b1)) || (rob_valids_2[6'h39] == 1'b0) : (((rob_branch_masks_2[6'h39] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h39] == 1'b1)) || (rob_valids_2[6'h39] == 1'b0)) &&
	  (ROBisOlder(6'h3a,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h3a] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h3a] == 1'b1)) || (rob_valids_2[6'h3a] == 1'b0) : (((rob_branch_masks_2[6'h3a] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h3a] == 1'b1)) || (rob_valids_2[6'h3a] == 1'b0)) &&
	  (ROBisOlder(6'h3b,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h3b] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h3b] == 1'b1)) || (rob_valids_2[6'h3b] == 1'b0) : (((rob_branch_masks_2[6'h3b] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h3b] == 1'b1)) || (rob_valids_2[6'h3b] == 1'b0)) &&
	  (ROBisOlder(6'h3c,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h3c] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h3c] == 1'b1)) || (rob_valids_2[6'h3c] == 1'b0) : (((rob_branch_masks_2[6'h3c] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h3c] == 1'b1)) || (rob_valids_2[6'h3c] == 1'b0)) &&
	  (ROBisOlder(6'h3d,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h3d] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h3d] == 1'b1)) || (rob_valids_2[6'h3d] == 1'b0) : (((rob_branch_masks_2[6'h3d] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h3d] == 1'b1)) || (rob_valids_2[6'h3d] == 1'b0)) &&
	  (ROBisOlder(6'h3e,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h3e] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h3e] == 1'b1)) || (rob_valids_2[6'h3e] == 1'b0) : (((rob_branch_masks_2[6'h3e] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h3e] == 1'b1)) || (rob_valids_2[6'h3e] == 1'b0)) &&
	  (ROBisOlder(6'h3f,soc2.core.rob.io_rob_tail_idx,root_id) ? (((rob_branch_masks_2[6'h3f] & root_br_mask) == root_br_mask) && (rob_valids_2[6'h3f] == 1'b1)) || (rob_valids_2[6'h3f] == 1'b0) : (((rob_branch_masks_2[6'h3f] & root_br_mask) != root_br_mask) && (rob_valids_2[6'h3f] == 1'b1)) || (rob_valids_2[6'h3f] == 1'b0)) &&
	  (soc1.core.rob.full && soc1.core.rob.rob_head_lsb == 1'b1 && soc1.core.rob.rob_tail_lsb == 1'b0 ? ((rob_branch_masks_1[soc1.core.rob.io_rob_tail_idx] & root_br_mask) == root_br_mask) && (rob_valids_1[soc1.core.rob.io_rob_tail_idx] == 1'b1) || (rob_valids_1[soc1.core.rob.io_rob_tail_idx] == 1'b0) : 1'b1) &&
	  (soc2.core.rob.full && soc2.core.rob.rob_head_lsb == 1'b1 && soc2.core.rob.rob_tail_lsb == 1'b0 ? ((rob_branch_masks_2[soc2.core.rob.io_rob_tail_idx] & root_br_mask) == root_br_mask) && (rob_valids_2[soc2.core.rob.io_rob_tail_idx] == 1'b1) || (rob_valids_2[soc2.core.rob.io_rob_tail_idx] == 1'b0) : 1'b1)
	  :
	  1'b1
	;

      //make sure that the branch at root_id commits only after its prediction is resolved as a misprediction
      wire root_commits_after_misprediction;
      assign root_commits_after_misprediction =
        (root_id[0] == 1'b0)
        ?
          (
          (soc1.core.rob.rob_head == root_id[5:1])
          ?
            soc1.core.rob.will_commit_0
            ?
              mispred_happened_1 == 1'b1
            :
              1'b1
          :
            1'b1
          ) &&
          (
          (soc2.core.rob.rob_head == root_id[5:1])
          ?
            soc2.core.rob.will_commit_0
            ?
              mispred_happened_2 == 1'b1
            :
              1'b1
          :
            1'b1
          )
        :
          (
          (soc1.core.rob.rob_head == root_id[5:1])
          ?
            soc1.core.rob.will_commit_1
            ?
              mispred_happened_1 == 1'b1
            :
              1'b1
          :
            1'b1
          ) &&
          (
          (soc2.core.rob.rob_head == root_id[5:1])
          ?
            soc2.core.rob.will_commit_1
            ?
              mispred_happened_2 == 1'b1
            :
              1'b1
          :
            1'b1
          )
      ;

      ///New stuff
      
	/*//check if a valid uop in ROB that uses STQ also exists in STQ
	function automatic ROB_exists_in_STQ(input [5:0] rob_idx, input rob_valids[63:0], input rob_uses_stq[63:0], input [1:0] rob_state, input _T_2387, input [5:0] stq_rob_idx[15:0], input [3:0] rob_stq_indexes[63:0], input stq_valids[15:0], input stq_committed[15:0]);
	begin
	  ROB_exists_in_STQ =
	  rob_valids[rob_idx] && rob_uses_stq[rob_idx] && rob_state != 2'h2 && _T_2387 != 1'b1
	  ?
	    stq_rob_idx[rob_stq_indexes[rob_idx]] == rob_idx && stq_valids[rob_stq_indexes[rob_idx]] && !stq_committed[rob_stq_indexes[rob_idx]]
	  :
	    1'b1
	  ;
	end
	endfunction

	//check if a valid uop in ROB that uses LDQ also exists in LDQ
	function automatic ROB_exists_in_LDQ(input [5:0] rob_idx, input rob_valids[63:0], input rob_uses_ldq[63:0], input [1:0] rob_state, input _T_2387, input rob_exception[63:0], input [5:0] ldq_rob_idx[15:0], input [3:0] rob_ldq_indexes[63:0], input ldq_valids[15:0]);
	begin
	  ROB_exists_in_LDQ =
	  rob_valids[rob_idx] && rob_uses_ldq[rob_idx] && rob_state != 2'h2 && _T_2387 != 1'b1 && !rob_exception[rob_idx]
	  ?
	    ldq_rob_idx[rob_ldq_indexes[rob_idx]] == rob_idx && ldq_valids[rob_ldq_indexes[rob_idx]]
	  :
	    1'b1
	  ;
	end
	endfunction*/

	//check if a valid uop in STQ also exists in ROB if not already committed
	function automatic STQ_exists_in_ROB(input [3:0] stq_idx, input stq_valids[15:0], input stq_committed[15:0], input rob_uses_stq[63:0], input [5:0] stq_rob_idx[15:0], input rob_valids[63:0]);
	begin
	  STQ_exists_in_ROB =
	  stq_valids[stq_idx] && !stq_committed[stq_idx]
	  ?
	    rob_uses_stq[stq_rob_idx[stq_idx]] && rob_valids[stq_rob_idx[stq_idx]]
	  :
	    1'b1
	  ;
	end
	endfunction

	//check if a valid uop in LDQ also exists in ROB if not already committed
	function automatic LDQ_exists_in_ROB(input [3:0] ldq_idx, input ldq_valids[15:0], input rob_uses_ldq[63:0], input [5:0] ldq_rob_idx[15:0], input rob_valids[63:0]);
	begin
	  LDQ_exists_in_ROB =
	  ldq_valids[ldq_idx]
	  ?
	    rob_uses_ldq[ldq_rob_idx[ldq_idx]] && rob_valids[ldq_rob_idx[ldq_idx]]
	  :
	    1'b1
	  ;
	end
	endfunction
	
	//check if a valid uop in a buffer also exists in ROB
	function automatic Buffer_exists_in_ROB(input buffer_valid, input buffer_uses_stq, input stq_committed[15:0], input [3:0] buffer_stq_idx, input rob_valids[63:0], input [5:0] buffer_rob_idx, 
	  input rob_uses_stq[63:0], input rob_uses_ldq[63:0], input buffer_uses_ldq);
	begin
	  Buffer_exists_in_ROB =
	  buffer_valid && !(buffer_uses_stq && stq_committed[buffer_stq_idx])
	  ?
	    rob_valids[buffer_rob_idx] &&
	    rob_uses_stq[buffer_rob_idx] == buffer_uses_stq &&
	    rob_uses_ldq[buffer_rob_idx] == buffer_uses_ldq
	  :
	    1'b1
	  ;
	end
	endfunction

	//check if a valid uop in a buffer also exists in ROB
	function automatic Buffer_exists_in_ROB_stq_idx_only(input buffer_valid, input stq_committed[15:0], input [3:0] buffer_stq_idx, input rob_valids[63:0], input [5:0] buffer_rob_idx);
	begin
	  Buffer_exists_in_ROB_stq_idx_only =
	  buffer_valid && !stq_committed[buffer_stq_idx]
	  ?
	    rob_valids[buffer_rob_idx]
	  :
	    1'b1
	  ;
	end
	endfunction

	//check if a valid uop in a buffer also exists in ROB
	function automatic Buffer_exists_in_ROB_only_uses_stq(input buffer_valid, input buffer_uses_stq, input rob_valids[63:0], input [5:0] buffer_rob_idx, input rob_uses_stq[63:0]);
	begin
	  Buffer_exists_in_ROB_only_uses_stq =
	  buffer_valid
	  ?
	    rob_valids[buffer_rob_idx] &&
	    rob_uses_stq[buffer_rob_idx] == buffer_uses_stq
	  :
	    1'b1
	  ;
	end
	endfunction

	//check if a valid uop in a buffer also exists in ROB
	function automatic Buffer_exists_in_ROB_only_stq(input buffer_valid, input buffer_uses_stq, input stq_committed[15:0], input [3:0] buffer_stq_idx, input rob_valids[63:0], input [5:0] buffer_rob_idx,
	  input rob_uses_stq[63:0]);
	begin
	  Buffer_exists_in_ROB_only_stq =
	  buffer_valid && !(buffer_uses_stq && stq_committed[buffer_stq_idx])
	  ?
	    rob_valids[buffer_rob_idx] &&
	    rob_uses_stq[buffer_rob_idx] == buffer_uses_stq
	  :
	    1'b1
	  ;
	end
	endfunction

	//check if a valid uop in a buffer also exists in ROB
	function automatic Buffer_exists_in_ROB_no_idx(input buffer_valid, input buffer_uses_stq, input rob_valids[63:0], input [5:0] buffer_rob_idx, input rob_uses_stq[63:0], input rob_uses_ldq[63:0], input buffer_uses_ldq);
	begin
	  Buffer_exists_in_ROB_no_idx =
	  buffer_valid
	  ?
	    rob_valids[buffer_rob_idx] &&
	    rob_uses_stq[buffer_rob_idx] == buffer_uses_stq &&
	    rob_uses_ldq[buffer_rob_idx] == buffer_uses_ldq
	  :
	    1'b1
	  ;
	end
	endfunction

	//check if a valid uop in a buffer also exists in LDQ
	function automatic Buffer_exists_in_LDQ(input buffer_valid, input buffer_uses_ldq, ldq_valids[15:0],  input [3:0] buffer_ldq_idx, ldq_uses_ldq[15:0]);
	begin
	  Buffer_exists_in_LDQ =
	  buffer_valid && buffer_uses_ldq
	  ?
	    ldq_valids[buffer_ldq_idx] &&
	    ldq_uses_ldq[buffer_ldq_idx]
	  :
	    1'b1
	  ;
	end
	endfunction

	//check if a valid uop in a buffer also exists in STQ
	function automatic Buffer_exists_in_STQ(input buffer_valid, input buffer_uses_stq, stq_valids[15:0],  input [3:0] buffer_stq_idx, stq_uses_stq[15:0]);
	begin
	  Buffer_exists_in_STQ =
	  buffer_valid && buffer_uses_stq
	  ?
	    stq_valids[buffer_stq_idx] &&
	    stq_uses_stq[buffer_stq_idx]
	  :
	    1'b1
	  ;
	end
	endfunction

        //Create an array of the branch masks of the ROB
	wire [11:0] rob_branch_masks_1 [63:0];
	assign rob_branch_masks_1[0] = soc1.core.rob.rob_uop__0_br_mask;
	assign rob_branch_masks_1[1] = soc1.core.rob.rob_uop_1_0_br_mask;
	assign rob_branch_masks_1[2] = soc1.core.rob.rob_uop__1_br_mask;
	assign rob_branch_masks_1[3] = soc1.core.rob.rob_uop_1_1_br_mask;
	assign rob_branch_masks_1[4] = soc1.core.rob.rob_uop__2_br_mask;
	assign rob_branch_masks_1[5] = soc1.core.rob.rob_uop_1_2_br_mask;
	assign rob_branch_masks_1[6] = soc1.core.rob.rob_uop__3_br_mask;
	assign rob_branch_masks_1[7] = soc1.core.rob.rob_uop_1_3_br_mask;
	assign rob_branch_masks_1[8] = soc1.core.rob.rob_uop__4_br_mask;
	assign rob_branch_masks_1[9] = soc1.core.rob.rob_uop_1_4_br_mask;
	assign rob_branch_masks_1[10] = soc1.core.rob.rob_uop__5_br_mask;
	assign rob_branch_masks_1[11] = soc1.core.rob.rob_uop_1_5_br_mask;
	assign rob_branch_masks_1[12] = soc1.core.rob.rob_uop__6_br_mask;
	assign rob_branch_masks_1[13] = soc1.core.rob.rob_uop_1_6_br_mask;
	assign rob_branch_masks_1[14] = soc1.core.rob.rob_uop__7_br_mask;
	assign rob_branch_masks_1[15] = soc1.core.rob.rob_uop_1_7_br_mask;
	assign rob_branch_masks_1[16] = soc1.core.rob.rob_uop__8_br_mask;
	assign rob_branch_masks_1[17] = soc1.core.rob.rob_uop_1_8_br_mask;
	assign rob_branch_masks_1[18] = soc1.core.rob.rob_uop__9_br_mask;
	assign rob_branch_masks_1[19] = soc1.core.rob.rob_uop_1_9_br_mask;
	assign rob_branch_masks_1[20] = soc1.core.rob.rob_uop__10_br_mask;
	assign rob_branch_masks_1[21] = soc1.core.rob.rob_uop_1_10_br_mask;
	assign rob_branch_masks_1[22] = soc1.core.rob.rob_uop__11_br_mask;
	assign rob_branch_masks_1[23] = soc1.core.rob.rob_uop_1_11_br_mask;
	assign rob_branch_masks_1[24] = soc1.core.rob.rob_uop__12_br_mask;
	assign rob_branch_masks_1[25] = soc1.core.rob.rob_uop_1_12_br_mask;
	assign rob_branch_masks_1[26] = soc1.core.rob.rob_uop__13_br_mask;
	assign rob_branch_masks_1[27] = soc1.core.rob.rob_uop_1_13_br_mask;
	assign rob_branch_masks_1[28] = soc1.core.rob.rob_uop__14_br_mask;
	assign rob_branch_masks_1[29] = soc1.core.rob.rob_uop_1_14_br_mask;
	assign rob_branch_masks_1[30] = soc1.core.rob.rob_uop__15_br_mask;
	assign rob_branch_masks_1[31] = soc1.core.rob.rob_uop_1_15_br_mask;
	assign rob_branch_masks_1[32] = soc1.core.rob.rob_uop__16_br_mask;
	assign rob_branch_masks_1[33] = soc1.core.rob.rob_uop_1_16_br_mask;
	assign rob_branch_masks_1[34] = soc1.core.rob.rob_uop__17_br_mask;
	assign rob_branch_masks_1[35] = soc1.core.rob.rob_uop_1_17_br_mask;
	assign rob_branch_masks_1[36] = soc1.core.rob.rob_uop__18_br_mask;
	assign rob_branch_masks_1[37] = soc1.core.rob.rob_uop_1_18_br_mask;
	assign rob_branch_masks_1[38] = soc1.core.rob.rob_uop__19_br_mask;
	assign rob_branch_masks_1[39] = soc1.core.rob.rob_uop_1_19_br_mask;
	assign rob_branch_masks_1[40] = soc1.core.rob.rob_uop__20_br_mask;
	assign rob_branch_masks_1[41] = soc1.core.rob.rob_uop_1_20_br_mask;
	assign rob_branch_masks_1[42] = soc1.core.rob.rob_uop__21_br_mask;
	assign rob_branch_masks_1[43] = soc1.core.rob.rob_uop_1_21_br_mask;
	assign rob_branch_masks_1[44] = soc1.core.rob.rob_uop__22_br_mask;
	assign rob_branch_masks_1[45] = soc1.core.rob.rob_uop_1_22_br_mask;
	assign rob_branch_masks_1[46] = soc1.core.rob.rob_uop__23_br_mask;
	assign rob_branch_masks_1[47] = soc1.core.rob.rob_uop_1_23_br_mask;
	assign rob_branch_masks_1[48] = soc1.core.rob.rob_uop__24_br_mask;
	assign rob_branch_masks_1[49] = soc1.core.rob.rob_uop_1_24_br_mask;
	assign rob_branch_masks_1[50] = soc1.core.rob.rob_uop__25_br_mask;
	assign rob_branch_masks_1[51] = soc1.core.rob.rob_uop_1_25_br_mask;
	assign rob_branch_masks_1[52] = soc1.core.rob.rob_uop__26_br_mask;
	assign rob_branch_masks_1[53] = soc1.core.rob.rob_uop_1_26_br_mask;
	assign rob_branch_masks_1[54] = soc1.core.rob.rob_uop__27_br_mask;
	assign rob_branch_masks_1[55] = soc1.core.rob.rob_uop_1_27_br_mask;
	assign rob_branch_masks_1[56] = soc1.core.rob.rob_uop__28_br_mask;
	assign rob_branch_masks_1[57] = soc1.core.rob.rob_uop_1_28_br_mask;
	assign rob_branch_masks_1[58] = soc1.core.rob.rob_uop__29_br_mask;
	assign rob_branch_masks_1[59] = soc1.core.rob.rob_uop_1_29_br_mask;
	assign rob_branch_masks_1[60] = soc1.core.rob.rob_uop__30_br_mask;
	assign rob_branch_masks_1[61] = soc1.core.rob.rob_uop_1_30_br_mask;
	assign rob_branch_masks_1[62] = soc1.core.rob.rob_uop__31_br_mask;
	assign rob_branch_masks_1[63] = soc1.core.rob.rob_uop_1_31_br_mask;

	//Create an array of the valid bits of the ROB
	wire rob_valids_1 [63:0];
	assign rob_valids_1[0] = soc1.core.rob.rob_val__0;
	assign rob_valids_1[1] = soc1.core.rob.rob_val_1_0;
	assign rob_valids_1[2] = soc1.core.rob.rob_val__1;
	assign rob_valids_1[3] = soc1.core.rob.rob_val_1_1;
	assign rob_valids_1[4] = soc1.core.rob.rob_val__2;
	assign rob_valids_1[5] = soc1.core.rob.rob_val_1_2;
	assign rob_valids_1[6] = soc1.core.rob.rob_val__3;
	assign rob_valids_1[7] = soc1.core.rob.rob_val_1_3;
	assign rob_valids_1[8] = soc1.core.rob.rob_val__4;
	assign rob_valids_1[9] = soc1.core.rob.rob_val_1_4;
	assign rob_valids_1[10] = soc1.core.rob.rob_val__5;
	assign rob_valids_1[11] = soc1.core.rob.rob_val_1_5;
	assign rob_valids_1[12] = soc1.core.rob.rob_val__6;
	assign rob_valids_1[13] = soc1.core.rob.rob_val_1_6;
	assign rob_valids_1[14] = soc1.core.rob.rob_val__7;
	assign rob_valids_1[15] = soc1.core.rob.rob_val_1_7;
	assign rob_valids_1[16] = soc1.core.rob.rob_val__8;
	assign rob_valids_1[17] = soc1.core.rob.rob_val_1_8;
	assign rob_valids_1[18] = soc1.core.rob.rob_val__9;
	assign rob_valids_1[19] = soc1.core.rob.rob_val_1_9;
	assign rob_valids_1[20] = soc1.core.rob.rob_val__10;
	assign rob_valids_1[21] = soc1.core.rob.rob_val_1_10;
	assign rob_valids_1[22] = soc1.core.rob.rob_val__11;
	assign rob_valids_1[23] = soc1.core.rob.rob_val_1_11;
	assign rob_valids_1[24] = soc1.core.rob.rob_val__12;
	assign rob_valids_1[25] = soc1.core.rob.rob_val_1_12;
	assign rob_valids_1[26] = soc1.core.rob.rob_val__13;
	assign rob_valids_1[27] = soc1.core.rob.rob_val_1_13;
	assign rob_valids_1[28] = soc1.core.rob.rob_val__14;
	assign rob_valids_1[29] = soc1.core.rob.rob_val_1_14;
	assign rob_valids_1[30] = soc1.core.rob.rob_val__15;
	assign rob_valids_1[31] = soc1.core.rob.rob_val_1_15;
	assign rob_valids_1[32] = soc1.core.rob.rob_val__16;
	assign rob_valids_1[33] = soc1.core.rob.rob_val_1_16;
	assign rob_valids_1[34] = soc1.core.rob.rob_val__17;
	assign rob_valids_1[35] = soc1.core.rob.rob_val_1_17;
	assign rob_valids_1[36] = soc1.core.rob.rob_val__18;
	assign rob_valids_1[37] = soc1.core.rob.rob_val_1_18;
	assign rob_valids_1[38] = soc1.core.rob.rob_val__19;
	assign rob_valids_1[39] = soc1.core.rob.rob_val_1_19;
	assign rob_valids_1[40] = soc1.core.rob.rob_val__20;
	assign rob_valids_1[41] = soc1.core.rob.rob_val_1_20;
	assign rob_valids_1[42] = soc1.core.rob.rob_val__21;
	assign rob_valids_1[43] = soc1.core.rob.rob_val_1_21;
	assign rob_valids_1[44] = soc1.core.rob.rob_val__22;
	assign rob_valids_1[45] = soc1.core.rob.rob_val_1_22;
	assign rob_valids_1[46] = soc1.core.rob.rob_val__23;
	assign rob_valids_1[47] = soc1.core.rob.rob_val_1_23;
	assign rob_valids_1[48] = soc1.core.rob.rob_val__24;
	assign rob_valids_1[49] = soc1.core.rob.rob_val_1_24;
	assign rob_valids_1[50] = soc1.core.rob.rob_val__25;
	assign rob_valids_1[51] = soc1.core.rob.rob_val_1_25;
	assign rob_valids_1[52] = soc1.core.rob.rob_val__26;
	assign rob_valids_1[53] = soc1.core.rob.rob_val_1_26;
	assign rob_valids_1[54] = soc1.core.rob.rob_val__27;
	assign rob_valids_1[55] = soc1.core.rob.rob_val_1_27;
	assign rob_valids_1[56] = soc1.core.rob.rob_val__28;
	assign rob_valids_1[57] = soc1.core.rob.rob_val_1_28;
	assign rob_valids_1[58] = soc1.core.rob.rob_val__29;
	assign rob_valids_1[59] = soc1.core.rob.rob_val_1_29;
	assign rob_valids_1[60] = soc1.core.rob.rob_val__30;
	assign rob_valids_1[61] = soc1.core.rob.rob_val_1_30;
	assign rob_valids_1[62] = soc1.core.rob.rob_val__31;
	assign rob_valids_1[63] = soc1.core.rob.rob_val_1_31;

	wire rob_uses_stq_1 [63:0];
	assign rob_uses_stq_1[0] = soc1.core.rob.rob_uop__0_uses_stq;
	assign rob_uses_stq_1[1] = soc1.core.rob.rob_uop_1_0_uses_stq;
	assign rob_uses_stq_1[2] = soc1.core.rob.rob_uop__1_uses_stq;
	assign rob_uses_stq_1[3] = soc1.core.rob.rob_uop_1_1_uses_stq;
	assign rob_uses_stq_1[4] = soc1.core.rob.rob_uop__2_uses_stq;
	assign rob_uses_stq_1[5] = soc1.core.rob.rob_uop_1_2_uses_stq;
	assign rob_uses_stq_1[6] = soc1.core.rob.rob_uop__3_uses_stq;
	assign rob_uses_stq_1[7] = soc1.core.rob.rob_uop_1_3_uses_stq;
	assign rob_uses_stq_1[8] = soc1.core.rob.rob_uop__4_uses_stq;
	assign rob_uses_stq_1[9] = soc1.core.rob.rob_uop_1_4_uses_stq;
	assign rob_uses_stq_1[10] = soc1.core.rob.rob_uop__5_uses_stq;
	assign rob_uses_stq_1[11] = soc1.core.rob.rob_uop_1_5_uses_stq;
	assign rob_uses_stq_1[12] = soc1.core.rob.rob_uop__6_uses_stq;
	assign rob_uses_stq_1[13] = soc1.core.rob.rob_uop_1_6_uses_stq;
	assign rob_uses_stq_1[14] = soc1.core.rob.rob_uop__7_uses_stq;
	assign rob_uses_stq_1[15] = soc1.core.rob.rob_uop_1_7_uses_stq;
	assign rob_uses_stq_1[16] = soc1.core.rob.rob_uop__8_uses_stq;
	assign rob_uses_stq_1[17] = soc1.core.rob.rob_uop_1_8_uses_stq;
	assign rob_uses_stq_1[18] = soc1.core.rob.rob_uop__9_uses_stq;
	assign rob_uses_stq_1[19] = soc1.core.rob.rob_uop_1_9_uses_stq;
	assign rob_uses_stq_1[20] = soc1.core.rob.rob_uop__10_uses_stq;
	assign rob_uses_stq_1[21] = soc1.core.rob.rob_uop_1_10_uses_stq;
	assign rob_uses_stq_1[22] = soc1.core.rob.rob_uop__11_uses_stq;
	assign rob_uses_stq_1[23] = soc1.core.rob.rob_uop_1_11_uses_stq;
	assign rob_uses_stq_1[24] = soc1.core.rob.rob_uop__12_uses_stq;
	assign rob_uses_stq_1[25] = soc1.core.rob.rob_uop_1_12_uses_stq;
	assign rob_uses_stq_1[26] = soc1.core.rob.rob_uop__13_uses_stq;
	assign rob_uses_stq_1[27] = soc1.core.rob.rob_uop_1_13_uses_stq;
	assign rob_uses_stq_1[28] = soc1.core.rob.rob_uop__14_uses_stq;
	assign rob_uses_stq_1[29] = soc1.core.rob.rob_uop_1_14_uses_stq;
	assign rob_uses_stq_1[30] = soc1.core.rob.rob_uop__15_uses_stq;
	assign rob_uses_stq_1[31] = soc1.core.rob.rob_uop_1_15_uses_stq;
	assign rob_uses_stq_1[32] = soc1.core.rob.rob_uop__16_uses_stq;
	assign rob_uses_stq_1[33] = soc1.core.rob.rob_uop_1_16_uses_stq;
	assign rob_uses_stq_1[34] = soc1.core.rob.rob_uop__17_uses_stq;
	assign rob_uses_stq_1[35] = soc1.core.rob.rob_uop_1_17_uses_stq;
	assign rob_uses_stq_1[36] = soc1.core.rob.rob_uop__18_uses_stq;
	assign rob_uses_stq_1[37] = soc1.core.rob.rob_uop_1_18_uses_stq;
	assign rob_uses_stq_1[38] = soc1.core.rob.rob_uop__19_uses_stq;
	assign rob_uses_stq_1[39] = soc1.core.rob.rob_uop_1_19_uses_stq;
	assign rob_uses_stq_1[40] = soc1.core.rob.rob_uop__20_uses_stq;
	assign rob_uses_stq_1[41] = soc1.core.rob.rob_uop_1_20_uses_stq;
	assign rob_uses_stq_1[42] = soc1.core.rob.rob_uop__21_uses_stq;
	assign rob_uses_stq_1[43] = soc1.core.rob.rob_uop_1_21_uses_stq;
	assign rob_uses_stq_1[44] = soc1.core.rob.rob_uop__22_uses_stq;
	assign rob_uses_stq_1[45] = soc1.core.rob.rob_uop_1_22_uses_stq;
	assign rob_uses_stq_1[46] = soc1.core.rob.rob_uop__23_uses_stq;
	assign rob_uses_stq_1[47] = soc1.core.rob.rob_uop_1_23_uses_stq;
	assign rob_uses_stq_1[48] = soc1.core.rob.rob_uop__24_uses_stq;
	assign rob_uses_stq_1[49] = soc1.core.rob.rob_uop_1_24_uses_stq;
	assign rob_uses_stq_1[50] = soc1.core.rob.rob_uop__25_uses_stq;
	assign rob_uses_stq_1[51] = soc1.core.rob.rob_uop_1_25_uses_stq;
	assign rob_uses_stq_1[52] = soc1.core.rob.rob_uop__26_uses_stq;
	assign rob_uses_stq_1[53] = soc1.core.rob.rob_uop_1_26_uses_stq;
	assign rob_uses_stq_1[54] = soc1.core.rob.rob_uop__27_uses_stq;
	assign rob_uses_stq_1[55] = soc1.core.rob.rob_uop_1_27_uses_stq;
	assign rob_uses_stq_1[56] = soc1.core.rob.rob_uop__28_uses_stq;
	assign rob_uses_stq_1[57] = soc1.core.rob.rob_uop_1_28_uses_stq;
	assign rob_uses_stq_1[58] = soc1.core.rob.rob_uop__29_uses_stq;
	assign rob_uses_stq_1[59] = soc1.core.rob.rob_uop_1_29_uses_stq;
	assign rob_uses_stq_1[60] = soc1.core.rob.rob_uop__30_uses_stq;
	assign rob_uses_stq_1[61] = soc1.core.rob.rob_uop_1_30_uses_stq;
	assign rob_uses_stq_1[62] = soc1.core.rob.rob_uop__31_uses_stq;
	assign rob_uses_stq_1[63] = soc1.core.rob.rob_uop_1_31_uses_stq;

	wire rob_uses_ldq_1 [63:0];
	assign rob_uses_ldq_1[0] = soc1.core.rob.rob_uop__0_uses_ldq;
	assign rob_uses_ldq_1[1] = soc1.core.rob.rob_uop_1_0_uses_ldq;
	assign rob_uses_ldq_1[2] = soc1.core.rob.rob_uop__1_uses_ldq;
	assign rob_uses_ldq_1[3] = soc1.core.rob.rob_uop_1_1_uses_ldq;
	assign rob_uses_ldq_1[4] = soc1.core.rob.rob_uop__2_uses_ldq;
	assign rob_uses_ldq_1[5] = soc1.core.rob.rob_uop_1_2_uses_ldq;
	assign rob_uses_ldq_1[6] = soc1.core.rob.rob_uop__3_uses_ldq;
	assign rob_uses_ldq_1[7] = soc1.core.rob.rob_uop_1_3_uses_ldq;
	assign rob_uses_ldq_1[8] = soc1.core.rob.rob_uop__4_uses_ldq;
	assign rob_uses_ldq_1[9] = soc1.core.rob.rob_uop_1_4_uses_ldq;
	assign rob_uses_ldq_1[10] = soc1.core.rob.rob_uop__5_uses_ldq;
	assign rob_uses_ldq_1[11] = soc1.core.rob.rob_uop_1_5_uses_ldq;
	assign rob_uses_ldq_1[12] = soc1.core.rob.rob_uop__6_uses_ldq;
	assign rob_uses_ldq_1[13] = soc1.core.rob.rob_uop_1_6_uses_ldq;
	assign rob_uses_ldq_1[14] = soc1.core.rob.rob_uop__7_uses_ldq;
	assign rob_uses_ldq_1[15] = soc1.core.rob.rob_uop_1_7_uses_ldq;
	assign rob_uses_ldq_1[16] = soc1.core.rob.rob_uop__8_uses_ldq;
	assign rob_uses_ldq_1[17] = soc1.core.rob.rob_uop_1_8_uses_ldq;
	assign rob_uses_ldq_1[18] = soc1.core.rob.rob_uop__9_uses_ldq;
	assign rob_uses_ldq_1[19] = soc1.core.rob.rob_uop_1_9_uses_ldq;
	assign rob_uses_ldq_1[20] = soc1.core.rob.rob_uop__10_uses_ldq;
	assign rob_uses_ldq_1[21] = soc1.core.rob.rob_uop_1_10_uses_ldq;
	assign rob_uses_ldq_1[22] = soc1.core.rob.rob_uop__11_uses_ldq;
	assign rob_uses_ldq_1[23] = soc1.core.rob.rob_uop_1_11_uses_ldq;
	assign rob_uses_ldq_1[24] = soc1.core.rob.rob_uop__12_uses_ldq;
	assign rob_uses_ldq_1[25] = soc1.core.rob.rob_uop_1_12_uses_ldq;
	assign rob_uses_ldq_1[26] = soc1.core.rob.rob_uop__13_uses_ldq;
	assign rob_uses_ldq_1[27] = soc1.core.rob.rob_uop_1_13_uses_ldq;
	assign rob_uses_ldq_1[28] = soc1.core.rob.rob_uop__14_uses_ldq;
	assign rob_uses_ldq_1[29] = soc1.core.rob.rob_uop_1_14_uses_ldq;
	assign rob_uses_ldq_1[30] = soc1.core.rob.rob_uop__15_uses_ldq;
	assign rob_uses_ldq_1[31] = soc1.core.rob.rob_uop_1_15_uses_ldq;
	assign rob_uses_ldq_1[32] = soc1.core.rob.rob_uop__16_uses_ldq;
	assign rob_uses_ldq_1[33] = soc1.core.rob.rob_uop_1_16_uses_ldq;
	assign rob_uses_ldq_1[34] = soc1.core.rob.rob_uop__17_uses_ldq;
	assign rob_uses_ldq_1[35] = soc1.core.rob.rob_uop_1_17_uses_ldq;
	assign rob_uses_ldq_1[36] = soc1.core.rob.rob_uop__18_uses_ldq;
	assign rob_uses_ldq_1[37] = soc1.core.rob.rob_uop_1_18_uses_ldq;
	assign rob_uses_ldq_1[38] = soc1.core.rob.rob_uop__19_uses_ldq;
	assign rob_uses_ldq_1[39] = soc1.core.rob.rob_uop_1_19_uses_ldq;
	assign rob_uses_ldq_1[40] = soc1.core.rob.rob_uop__20_uses_ldq;
	assign rob_uses_ldq_1[41] = soc1.core.rob.rob_uop_1_20_uses_ldq;
	assign rob_uses_ldq_1[42] = soc1.core.rob.rob_uop__21_uses_ldq;
	assign rob_uses_ldq_1[43] = soc1.core.rob.rob_uop_1_21_uses_ldq;
	assign rob_uses_ldq_1[44] = soc1.core.rob.rob_uop__22_uses_ldq;
	assign rob_uses_ldq_1[45] = soc1.core.rob.rob_uop_1_22_uses_ldq;
	assign rob_uses_ldq_1[46] = soc1.core.rob.rob_uop__23_uses_ldq;
	assign rob_uses_ldq_1[47] = soc1.core.rob.rob_uop_1_23_uses_ldq;
	assign rob_uses_ldq_1[48] = soc1.core.rob.rob_uop__24_uses_ldq;
	assign rob_uses_ldq_1[49] = soc1.core.rob.rob_uop_1_24_uses_ldq;
	assign rob_uses_ldq_1[50] = soc1.core.rob.rob_uop__25_uses_ldq;
	assign rob_uses_ldq_1[51] = soc1.core.rob.rob_uop_1_25_uses_ldq;
	assign rob_uses_ldq_1[52] = soc1.core.rob.rob_uop__26_uses_ldq;
	assign rob_uses_ldq_1[53] = soc1.core.rob.rob_uop_1_26_uses_ldq;
	assign rob_uses_ldq_1[54] = soc1.core.rob.rob_uop__27_uses_ldq;
	assign rob_uses_ldq_1[55] = soc1.core.rob.rob_uop_1_27_uses_ldq;
	assign rob_uses_ldq_1[56] = soc1.core.rob.rob_uop__28_uses_ldq;
	assign rob_uses_ldq_1[57] = soc1.core.rob.rob_uop_1_28_uses_ldq;
	assign rob_uses_ldq_1[58] = soc1.core.rob.rob_uop__29_uses_ldq;
	assign rob_uses_ldq_1[59] = soc1.core.rob.rob_uop_1_29_uses_ldq;
	assign rob_uses_ldq_1[60] = soc1.core.rob.rob_uop__30_uses_ldq;
	assign rob_uses_ldq_1[61] = soc1.core.rob.rob_uop_1_30_uses_ldq;
	assign rob_uses_ldq_1[62] = soc1.core.rob.rob_uop__31_uses_ldq;
	assign rob_uses_ldq_1[63] = soc1.core.rob.rob_uop_1_31_uses_ldq;
	
	//Create an array of the exception bits of the ROB
	wire rob_exception_1 [63:0];
	assign rob_exception_1[0] = soc1.core.rob.rob_exception__0;
	assign rob_exception_1[1] = soc1.core.rob.rob_exception_1_0;
	assign rob_exception_1[2] = soc1.core.rob.rob_exception__1;
	assign rob_exception_1[3] = soc1.core.rob.rob_exception_1_1;
	assign rob_exception_1[4] = soc1.core.rob.rob_exception__2;
	assign rob_exception_1[5] = soc1.core.rob.rob_exception_1_2;
	assign rob_exception_1[6] = soc1.core.rob.rob_exception__3;
	assign rob_exception_1[7] = soc1.core.rob.rob_exception_1_3;
	assign rob_exception_1[8] = soc1.core.rob.rob_exception__4;
	assign rob_exception_1[9] = soc1.core.rob.rob_exception_1_4;
	assign rob_exception_1[10] = soc1.core.rob.rob_exception__5;
	assign rob_exception_1[11] = soc1.core.rob.rob_exception_1_5;
	assign rob_exception_1[12] = soc1.core.rob.rob_exception__6;
	assign rob_exception_1[13] = soc1.core.rob.rob_exception_1_6;
	assign rob_exception_1[14] = soc1.core.rob.rob_exception__7;
	assign rob_exception_1[15] = soc1.core.rob.rob_exception_1_7;
	assign rob_exception_1[16] = soc1.core.rob.rob_exception__8;
	assign rob_exception_1[17] = soc1.core.rob.rob_exception_1_8;
	assign rob_exception_1[18] = soc1.core.rob.rob_exception__9;
	assign rob_exception_1[19] = soc1.core.rob.rob_exception_1_9;
	assign rob_exception_1[20] = soc1.core.rob.rob_exception__10;
	assign rob_exception_1[21] = soc1.core.rob.rob_exception_1_10;
	assign rob_exception_1[22] = soc1.core.rob.rob_exception__11;
	assign rob_exception_1[23] = soc1.core.rob.rob_exception_1_11;
	assign rob_exception_1[24] = soc1.core.rob.rob_exception__12;
	assign rob_exception_1[25] = soc1.core.rob.rob_exception_1_12;
	assign rob_exception_1[26] = soc1.core.rob.rob_exception__13;
	assign rob_exception_1[27] = soc1.core.rob.rob_exception_1_13;
	assign rob_exception_1[28] = soc1.core.rob.rob_exception__14;
	assign rob_exception_1[29] = soc1.core.rob.rob_exception_1_14;
	assign rob_exception_1[30] = soc1.core.rob.rob_exception__15;
	assign rob_exception_1[31] = soc1.core.rob.rob_exception_1_15;
	assign rob_exception_1[32] = soc1.core.rob.rob_exception__16;
	assign rob_exception_1[33] = soc1.core.rob.rob_exception_1_16;
	assign rob_exception_1[34] = soc1.core.rob.rob_exception__17;
	assign rob_exception_1[35] = soc1.core.rob.rob_exception_1_17;
	assign rob_exception_1[36] = soc1.core.rob.rob_exception__18;
	assign rob_exception_1[37] = soc1.core.rob.rob_exception_1_18;
	assign rob_exception_1[38] = soc1.core.rob.rob_exception__19;
	assign rob_exception_1[39] = soc1.core.rob.rob_exception_1_19;
	assign rob_exception_1[40] = soc1.core.rob.rob_exception__20;
	assign rob_exception_1[41] = soc1.core.rob.rob_exception_1_20;
	assign rob_exception_1[42] = soc1.core.rob.rob_exception__21;
	assign rob_exception_1[43] = soc1.core.rob.rob_exception_1_21;
	assign rob_exception_1[44] = soc1.core.rob.rob_exception__22;
	assign rob_exception_1[45] = soc1.core.rob.rob_exception_1_22;
	assign rob_exception_1[46] = soc1.core.rob.rob_exception__23;
	assign rob_exception_1[47] = soc1.core.rob.rob_exception_1_23;
	assign rob_exception_1[48] = soc1.core.rob.rob_exception__24;
	assign rob_exception_1[49] = soc1.core.rob.rob_exception_1_24;
	assign rob_exception_1[50] = soc1.core.rob.rob_exception__25;
	assign rob_exception_1[51] = soc1.core.rob.rob_exception_1_25;
	assign rob_exception_1[52] = soc1.core.rob.rob_exception__26;
	assign rob_exception_1[53] = soc1.core.rob.rob_exception_1_26;
	assign rob_exception_1[54] = soc1.core.rob.rob_exception__27;
	assign rob_exception_1[55] = soc1.core.rob.rob_exception_1_27;
	assign rob_exception_1[56] = soc1.core.rob.rob_exception__28;
	assign rob_exception_1[57] = soc1.core.rob.rob_exception_1_28;
	assign rob_exception_1[58] = soc1.core.rob.rob_exception__29;
	assign rob_exception_1[59] = soc1.core.rob.rob_exception_1_29;
	assign rob_exception_1[60] = soc1.core.rob.rob_exception__30;
	assign rob_exception_1[61] = soc1.core.rob.rob_exception_1_30;
	assign rob_exception_1[62] = soc1.core.rob.rob_exception__31;
	assign rob_exception_1[63] = soc1.core.rob.rob_exception_1_31;

	//array that stores a copy of the rob_idx of the ldq
	wire [5:0] ldq_rob_idx_1 [15:0];
	assign ldq_rob_idx_1[0] = soc1.lsu.ldq_0_bits_uop_rob_idx;
	assign ldq_rob_idx_1[1] = soc1.lsu.ldq_1_bits_uop_rob_idx;
	assign ldq_rob_idx_1[2] = soc1.lsu.ldq_2_bits_uop_rob_idx;
	assign ldq_rob_idx_1[3] = soc1.lsu.ldq_3_bits_uop_rob_idx;
	assign ldq_rob_idx_1[4] = soc1.lsu.ldq_4_bits_uop_rob_idx;
	assign ldq_rob_idx_1[5] = soc1.lsu.ldq_5_bits_uop_rob_idx;
	assign ldq_rob_idx_1[6] = soc1.lsu.ldq_6_bits_uop_rob_idx;
	assign ldq_rob_idx_1[7] = soc1.lsu.ldq_7_bits_uop_rob_idx;
	assign ldq_rob_idx_1[8] = soc1.lsu.ldq_8_bits_uop_rob_idx;
	assign ldq_rob_idx_1[9] = soc1.lsu.ldq_9_bits_uop_rob_idx;
	assign ldq_rob_idx_1[10] = soc1.lsu.ldq_10_bits_uop_rob_idx;
	assign ldq_rob_idx_1[11] = soc1.lsu.ldq_11_bits_uop_rob_idx;
	assign ldq_rob_idx_1[12] = soc1.lsu.ldq_12_bits_uop_rob_idx;
	assign ldq_rob_idx_1[13] = soc1.lsu.ldq_13_bits_uop_rob_idx;
	assign ldq_rob_idx_1[14] = soc1.lsu.ldq_14_bits_uop_rob_idx;
	assign ldq_rob_idx_1[15] = soc1.lsu.ldq_15_bits_uop_rob_idx;

	//array that stores a copy of the rob_idx of the stq
	wire [5:0] stq_rob_idx_1 [15:0];
	assign stq_rob_idx_1[0] = soc1.lsu.stq_0_bits_uop_rob_idx;
	assign stq_rob_idx_1[1] = soc1.lsu.stq_1_bits_uop_rob_idx;
	assign stq_rob_idx_1[2] = soc1.lsu.stq_2_bits_uop_rob_idx;
	assign stq_rob_idx_1[3] = soc1.lsu.stq_3_bits_uop_rob_idx;
	assign stq_rob_idx_1[4] = soc1.lsu.stq_4_bits_uop_rob_idx;
	assign stq_rob_idx_1[5] = soc1.lsu.stq_5_bits_uop_rob_idx;
	assign stq_rob_idx_1[6] = soc1.lsu.stq_6_bits_uop_rob_idx;
	assign stq_rob_idx_1[7] = soc1.lsu.stq_7_bits_uop_rob_idx;
	assign stq_rob_idx_1[8] = soc1.lsu.stq_8_bits_uop_rob_idx;
	assign stq_rob_idx_1[9] = soc1.lsu.stq_9_bits_uop_rob_idx;
	assign stq_rob_idx_1[10] = soc1.lsu.stq_10_bits_uop_rob_idx;
	assign stq_rob_idx_1[11] = soc1.lsu.stq_11_bits_uop_rob_idx;
	assign stq_rob_idx_1[12] = soc1.lsu.stq_12_bits_uop_rob_idx;
	assign stq_rob_idx_1[13] = soc1.lsu.stq_13_bits_uop_rob_idx;
	assign stq_rob_idx_1[14] = soc1.lsu.stq_14_bits_uop_rob_idx;
	assign stq_rob_idx_1[15] = soc1.lsu.stq_15_bits_uop_rob_idx;

	//array that stores a copy of the committed bits of the stq
	wire stq_committed_1 [15:0];
	assign stq_committed_1[0] = soc1.lsu.stq_0_bits_committed;
	assign stq_committed_1[1] = soc1.lsu.stq_1_bits_committed;
	assign stq_committed_1[2] = soc1.lsu.stq_2_bits_committed;
	assign stq_committed_1[3] = soc1.lsu.stq_3_bits_committed;
	assign stq_committed_1[4] = soc1.lsu.stq_4_bits_committed;
	assign stq_committed_1[5] = soc1.lsu.stq_5_bits_committed;
	assign stq_committed_1[6] = soc1.lsu.stq_6_bits_committed;
	assign stq_committed_1[7] = soc1.lsu.stq_7_bits_committed;
	assign stq_committed_1[8] = soc1.lsu.stq_8_bits_committed;
	assign stq_committed_1[9] = soc1.lsu.stq_9_bits_committed;
	assign stq_committed_1[10] = soc1.lsu.stq_10_bits_committed;
	assign stq_committed_1[11] = soc1.lsu.stq_11_bits_committed;
	assign stq_committed_1[12] = soc1.lsu.stq_12_bits_committed;
	assign stq_committed_1[13] = soc1.lsu.stq_13_bits_committed;
	assign stq_committed_1[14] = soc1.lsu.stq_14_bits_committed;
	assign stq_committed_1[15] = soc1.lsu.stq_15_bits_committed;

	//function that returns true if the given ID in ROB is above or equal ldq_head and below ldq_tail
	function automatic isInBoundsROB_1;
	  //6-bit ID of the ROB entry
	  input [5:0] id;
	  begin
	    if(rob_valids_1[id] == 1'b1)
	    begin
	      //distinguish between positions of head and tail
	      if (soc1.core.rob.io_rob_head_idx < soc1.core.rob.io_rob_tail_idx)
	      begin
	  isInBoundsROB_1 = (id >= soc1.core.rob.io_rob_head_idx && id < soc1.core.rob.io_rob_tail_idx) || soc1.core.rob.full;
	      end
	      else if (soc1.core.rob.io_rob_head_idx > soc1.core.rob.io_rob_tail_idx)
	      begin
	  isInBoundsROB_1 = (id >= soc1.core.rob.io_rob_head_idx || id < soc1.core.rob.io_rob_tail_idx) || soc1.core.rob.full;
	      end
	      else // soc1.core.rob.io_rob_head_idx == soc1.core.rob.io_rob_tail_idx
	      begin
	  isInBoundsROB_1 = !soc1.core.rob.io_empty;
	      end
	    end
	    else
	    begin
	      isInBoundsROB_1 = 1'b0;
	    end
	  end
	endfunction

	function automatic ROBisOlder(input [5:0] id1, id2, head);
	begin
	  ROBisOlder = ((id1 < id2) ^ (id1 < head) ^ (id2 < head));
	end
	endfunction

  wire consistent_branch_masks_1;
	assign consistent_branch_masks_1 =
	(
	//is the uop at head valid and is the ROB not empty
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 0) % 64)
	?
	  (
	  //if true, the branch mask at head must be 0 because the first valid instruction after head must be non-speculative
	  rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 0) % 64] == 12'b0
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 1) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 0) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 0) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 1) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 0) % 64]
	  :
	    (
	    //if head is invalid, the branch mask at head + 1 must be 0 because the first valid instruction after head must be non-speculative
	    rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] == 12'b0
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 2) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 2) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 1) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 0) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 0) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 2) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 0) % 64]
	    :
	      //if head is invalid, the branch mask at head + 2 must be 0 because the first valid instruction after head must be non-speculative
	      rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] == 12'b0
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 3) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 3) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 2) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 3) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 1) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 0) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 3) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 0) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 4) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 4) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 3) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 4) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 2) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 4) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 1) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 5) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 5) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 4) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 5) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 3) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 5) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 2) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 6) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 6) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 5) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 6) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 4) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 6) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 3) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 7) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 7) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 6) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 7) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 5) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 7) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 4) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 8) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 8) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 7) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 8) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 6) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 8) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 5) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 9) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 9) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 8) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 9) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 7) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 9) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 6) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 10) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 10) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 9) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 10) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 8) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 10) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 7) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 11) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 11) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 10) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 11) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 9) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 11) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 8) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 12) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 12) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 11) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 12) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 10) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 12) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 9) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 13) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 13) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 12) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 13) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 11) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 13) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 10) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 14) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 14) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 13) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 14) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 12) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 14) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 11) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 15) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 15) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 14) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 15) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 13) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 15) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 12) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 16) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 16) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 15) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 16) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 14) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 16) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 13) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 17) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 17) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 16) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 17) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 15) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 17) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 14) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 18) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 18) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 17) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 18) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 16) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 18) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 15) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 19) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 19) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 18) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 19) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 17) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 19) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 16) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 20) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 20) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 19) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 20) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 18) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 20) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 17) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 21) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 21) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 20) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 21) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 19) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 21) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 18) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 22) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 22) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 21) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 22) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 20) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 22) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 19) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 23) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 23) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 22) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 23) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 21) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 23) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 20) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 24) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 24) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 23) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 24) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 22) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 24) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 21) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 25) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 25) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 24) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 25) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 23) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 25) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 22) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 26) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 26) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 25) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 26) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 24) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 26) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 23) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 27) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 27) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 26) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 27) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 25) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 27) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 24) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 28) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 28) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 27) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 28) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 26) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 28) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 25) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 29) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 29) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 28) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 29) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 27) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 29) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 26) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 30) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 30) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 29) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 30) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 28) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 30) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 27) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 31) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 31) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 30) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 31) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 29) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 31) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 28) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 32) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 32) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 31) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 32) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 30) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 32) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 29) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 33) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 33) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 32) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 33) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 31) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 33) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 30) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 34) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 34) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 33) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 34) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 32) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 34) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 31) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 35) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 35) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 34) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 35) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 33) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 35) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 32) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 36) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 36) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 35) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 36) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 34) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 36) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 33) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 37) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 37) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 36) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 37) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 35) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 37) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 34) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 38) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 38) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 37) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 38) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 36) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 38) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 35) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 39) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 39) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 38) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 39) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 37) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 39) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 36) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 40) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 40) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 39) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 40) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 38) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 40) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 37) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 41) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 41) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 40) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 41) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 39) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 41) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 38) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 42) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 42) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 41) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 42) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 40) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 42) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 39) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 43) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 43) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 42) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 43) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 41) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 43) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 40) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 44) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 44) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 43) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 44) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 42) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 44) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 41) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 45) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 45) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 44) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 45) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 43) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 45) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 42) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 46) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 46) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 45) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 46) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 44) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 46) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 43) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 47) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 47) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 46) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 47) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 45) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 47) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 44) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 48) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 48) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 47) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 48) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 46) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 48) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 45) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 49) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 49) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 48) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 49) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 47) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 49) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 46) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 50) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 50) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 49) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 50) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 48) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 50) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 47) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 51) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 51) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 50) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 51) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 49) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 51) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 48) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 52) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 52) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 51) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 52) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 50) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 52) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 49) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 53) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 53) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 52) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 53) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 51) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 53) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 50) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 54) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 54) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 53) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 54) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 52) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 54) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 51) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 55) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 55) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 54) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 55) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 53) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 55) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 52) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 56) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 56) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 55) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 56) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 54) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 56) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 53) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 57) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 57) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 56) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 57) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 55) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 57) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 54) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 58) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 58) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 57) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 58) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 56) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 58) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 55) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 59) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 59) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 58) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 59) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 57) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 59) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 56) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 60) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 60) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 59) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 60) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 58) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 60) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 57) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 61) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 61) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 60) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 61) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 59) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 61) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 58) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 62) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 61) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 62) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 61) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 62) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 60) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 62) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 59) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_1((soc1.core.rob.io_rob_head_idx + 63) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_1[(soc1.core.rob.io_rob_head_idx + 62) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 62) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 63) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 62) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 61) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 63) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 61) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] & rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 63) % 64]) == rob_branch_masks_1[(soc1.core.rob.io_rob_head_idx + 60) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	);

	wire consistent_valid_flags_1;
	assign consistent_valid_flags_1 =
	(
	soc1.core.rob.io_empty == 1'b1
	?
		//if empty, no entry can be valid
		(soc1.core.rob.rob_val__0 | soc1.core.rob.rob_val_1_0 | soc1.core.rob.rob_val__1 | soc1.core.rob.rob_val_1_1 | soc1.core.rob.rob_val__2 | soc1.core.rob.rob_val_1_2 |
		soc1.core.rob.rob_val__3 | soc1.core.rob.rob_val_1_3 | soc1.core.rob.rob_val__4 | soc1.core.rob.rob_val_1_4 | soc1.core.rob.rob_val__5 | soc1.core.rob.rob_val_1_5 |
		soc1.core.rob.rob_val__6 | soc1.core.rob.rob_val_1_6 | soc1.core.rob.rob_val__7 | soc1.core.rob.rob_val_1_7 | soc1.core.rob.rob_val__8 | soc1.core.rob.rob_val_1_8 |
		soc1.core.rob.rob_val__9 | soc1.core.rob.rob_val_1_9 | soc1.core.rob.rob_val__10 | soc1.core.rob.rob_val_1_10 | soc1.core.rob.rob_val__11 | soc1.core.rob.rob_val_1_11 |
		soc1.core.rob.rob_val__12 | soc1.core.rob.rob_val_1_12 | soc1.core.rob.rob_val__13 | soc1.core.rob.rob_val_1_13 | soc1.core.rob.rob_val__14 | soc1.core.rob.rob_val_1_14 |
		soc1.core.rob.rob_val__15 | soc1.core.rob.rob_val_1_15 | soc1.core.rob.rob_val__16 | soc1.core.rob.rob_val_1_16 | soc1.core.rob.rob_val__17 | soc1.core.rob.rob_val_1_17 |
		soc1.core.rob.rob_val__18 | soc1.core.rob.rob_val_1_18 | soc1.core.rob.rob_val__19 | soc1.core.rob.rob_val_1_19 | soc1.core.rob.rob_val__20 | soc1.core.rob.rob_val_1_20 |
		soc1.core.rob.rob_val__21 | soc1.core.rob.rob_val_1_21 | soc1.core.rob.rob_val__22 | soc1.core.rob.rob_val_1_22 | soc1.core.rob.rob_val__23 | soc1.core.rob.rob_val_1_23 |
		soc1.core.rob.rob_val__24 | soc1.core.rob.rob_val_1_24 | soc1.core.rob.rob_val__25 | soc1.core.rob.rob_val_1_25 | soc1.core.rob.rob_val__26 | soc1.core.rob.rob_val_1_26 |
		soc1.core.rob.rob_val__27 | soc1.core.rob.rob_val_1_27 | soc1.core.rob.rob_val__28 | soc1.core.rob.rob_val_1_28 | soc1.core.rob.rob_val__29 | soc1.core.rob.rob_val_1_29 |
		soc1.core.rob.rob_val__30 | soc1.core.rob.rob_val_1_30 | soc1.core.rob.rob_val__31 | soc1.core.rob.rob_val_1_31) == 1'b0
	:
		//if not empty
		//check for branch misprediction
		soc1.core.b2_mispredict
		?
			//only entries that are older than the mispredicted branch and the mispredicted branch itself can be valid
			//distinction for different head_lsbs
			(soc1.core.rob.rob_head_lsb == 1'b0)
			?
				//if not empty, at least one entry at head is valid
				//check for every entry if it is older than b2_uop_rob_idx + 1
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 0) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 0) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 0) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 1) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 0) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 1) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 2) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 2) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 4) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 4) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 6) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 6) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 8) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 8) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 10) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 10) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 12) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 12) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 14) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 14) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 16) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 16) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 18) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 18) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 20) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 20) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 22) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 22) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 24) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 24) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 26) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 26) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 28) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 28) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 30) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 30) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 32) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 32) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 34) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 34) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 36) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 36) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 38) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 38) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 40) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 40) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 42) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 42) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 44) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 44) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 46) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 46) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 48) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 48) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 50) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 50) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 52) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 52) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 54) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 54) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 56) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 56) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 58) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 58) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 60) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 60) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 62) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 62) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 62) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 63) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 62) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 63) % 64])
				)
			:
				//else if rob_head_lsb==1'b1
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 0) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 0) % 64) == soc1.core.b2_uop_rob_idx
				? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 0) % 64]
				: !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 0) % 64]
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 1) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 1) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 3) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 3) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 5) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 5) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 7) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 7) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 9) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 9) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 11) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 11) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 13) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 13) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 15) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 15) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 17) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 17) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 19) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 19) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 21) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 21) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 23) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 23) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 25) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 25) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 27) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 27) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 29) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 29) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 31) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 31) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 33) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 33) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 35) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 35) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 37) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 37) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 39) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 39) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 41) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 41) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 43) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 43) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 45) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 45) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 47) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 47) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 49) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 49) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 51) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 51) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 53) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 53) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 55) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 55) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 57) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 57) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 59) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 59) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 61) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 61) % 64) == soc1.core.b2_uop_rob_idx
				? (rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 62) % 64])
				: (!rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 62) % 64])
				) &&
				(ROBisOlder((soc1.core.rob.io_rob_head_idx + 63) % 64, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) || ((soc1.core.rob.io_rob_head_idx + 63) % 64) == soc1.core.b2_uop_rob_idx
				? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 63) % 64]
				: !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 63) % 64]
				)
		:
			soc1.core.rob.full == 1'b1
			?
				//if full, at least one entry per row has to be valid
				(soc1.core.rob.rob_val__0 || soc1.core.rob.rob_val_1_0) && (soc1.core.rob.rob_val__1 || soc1.core.rob.rob_val_1_1) && (soc1.core.rob.rob_val__2 || soc1.core.rob.rob_val_1_2) &&
				(soc1.core.rob.rob_val__3 || soc1.core.rob.rob_val_1_3) && (soc1.core.rob.rob_val__4 || soc1.core.rob.rob_val_1_4) && (soc1.core.rob.rob_val__5 || soc1.core.rob.rob_val_1_5) &&
				(soc1.core.rob.rob_val__6 || soc1.core.rob.rob_val_1_6) && (soc1.core.rob.rob_val__7 || soc1.core.rob.rob_val_1_7) && (soc1.core.rob.rob_val__8 || soc1.core.rob.rob_val_1_8) &&
				(soc1.core.rob.rob_val__9 || soc1.core.rob.rob_val_1_9) && (soc1.core.rob.rob_val__10 || soc1.core.rob.rob_val_1_10) && (soc1.core.rob.rob_val__11 || soc1.core.rob.rob_val_1_11) &&
				(soc1.core.rob.rob_val__12 || soc1.core.rob.rob_val_1_12) && (soc1.core.rob.rob_val__13 || soc1.core.rob.rob_val_1_13) && (soc1.core.rob.rob_val__14 || soc1.core.rob.rob_val_1_14) &&
				(soc1.core.rob.rob_val__15 || soc1.core.rob.rob_val_1_15) && (soc1.core.rob.rob_val__16 || soc1.core.rob.rob_val_1_16) && (soc1.core.rob.rob_val__17 || soc1.core.rob.rob_val_1_17) &&
				(soc1.core.rob.rob_val__18 || soc1.core.rob.rob_val_1_18) && (soc1.core.rob.rob_val__19 || soc1.core.rob.rob_val_1_19) && (soc1.core.rob.rob_val__20 || soc1.core.rob.rob_val_1_20) &&
				(soc1.core.rob.rob_val__21 || soc1.core.rob.rob_val_1_21) && (soc1.core.rob.rob_val__22 || soc1.core.rob.rob_val_1_22) && (soc1.core.rob.rob_val__23 || soc1.core.rob.rob_val_1_23) &&
				(soc1.core.rob.rob_val__24 || soc1.core.rob.rob_val_1_24) && (soc1.core.rob.rob_val__25 || soc1.core.rob.rob_val_1_25) && (soc1.core.rob.rob_val__26 || soc1.core.rob.rob_val_1_26) &&
				(soc1.core.rob.rob_val__27 || soc1.core.rob.rob_val_1_27) && (soc1.core.rob.rob_val__28 || soc1.core.rob.rob_val_1_28) && (soc1.core.rob.rob_val__29 || soc1.core.rob.rob_val_1_29) &&
				(soc1.core.rob.rob_val__30 || soc1.core.rob.rob_val_1_30) && (soc1.core.rob.rob_val__31 || soc1.core.rob.rob_val_1_31)
			:
				//if not empty, full, rollback or branch mispredict
				//in every row, that is older than tail there has to be at least one valid entry
				//distinction for different head_lsbs
				(
				(soc1.core.rob.rob_head_lsb == 1'b0)
				?
					//if neither full or empty, at least one entry at head is valid
					(rob_valids_1[(soc1.core.rob.io_rob_head_idx + 0) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 1) % 64]) &&
					//for every row that is before tail, there is at least one valid entry
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 2) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 4) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 6) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 8) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 10) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 12) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 14) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 16) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 18) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 20) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 22) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 24) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 26) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 28) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 30) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 32) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 34) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 36) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 38) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 40) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 42) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 44) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 46) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 48) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 50) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 52) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 54) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 56) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 58) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 60) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 62) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 62) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 63) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 62) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 63) % 64]) &&
					//make sure that tail points an invalid entry
					(soc1.core.rob.rob_state == 2'h2 ? 1'b1 : rob_valids_1[soc1.core.rob.io_rob_tail_idx] == 1'b0)
				:
					//if soc1.core.rob.rob_head_lsb == 1'b1
					//if neither full or empty, head must be valid, since head_lsb is 1
					(rob_valids_1[(soc1.core.rob.io_rob_head_idx + 0) % 64]) &&
					//for every row that is before tail, there is at least one valid entry
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 1) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 1) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 2) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 3) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 3) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 4) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 5) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 5) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 6) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 7) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 7) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 8) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 9) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 9) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 10) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 11) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 11) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 12) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 13) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 13) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 14) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 15) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 15) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 16) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 17) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 17) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 18) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 19) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 19) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 20) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 21) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 21) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 22) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 23) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 23) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 24) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 25) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 25) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 26) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 27) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 27) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 28) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 29) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 29) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 30) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 31) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 31) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 32) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 33) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 33) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 34) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 35) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 35) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 36) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 37) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 37) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 38) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 39) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 39) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 40) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 41) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 41) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 42) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 43) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 43) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 44) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 45) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 45) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 46) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 47) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 47) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 48) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 49) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 49) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 50) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 51) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 51) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 52) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 53) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 53) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 54) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 55) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 55) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 56) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 57) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 57) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 58) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 59) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 59) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 60) % 64]) &&
					((ROBisOlder((soc1.core.rob.io_rob_head_idx + 61) % 64, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx)) ? rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64] || rob_valids_1[(soc1.core.rob.io_rob_head_idx + 62) % 64] : !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 61) % 64] && !rob_valids_1[(soc1.core.rob.io_rob_head_idx + 62) % 64]) &&
					//head+63 is in fact the entry before head+0, which must be invalid, since ROB is not full
					(rob_valids_1[(soc1.core.rob.io_rob_head_idx + 63) % 64] == 1'b0) &&
					//make sure that tail points an invalid entry
					(soc1.core.rob.rob_state == 2'h2 ? 1'b1 : rob_valids_1[soc1.core.rob.io_rob_tail_idx] == 1'b0)
				)
	);


	//if tail is rolled back because of a mispredict, make sure it is rolled back to an older value than tail
	wire consistent_tail_rollback_1;
	assign consistent_tail_rollback_1 =
	  (soc1.core.b2_mispredict == 1'b1 ? ROBisOlder(soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx) || soc1.core.rob.full: 1'b1)
	;

	//ensure that no speculative instruction commits
	wire no_speculative_commit_1;
	assign no_speculative_commit_1 =
	  (soc1.core.rob.will_commit_0 ? (rob_branch_masks_1[{soc1.core.rob.rob_head, 1'b0}] == 12'b0) && rob_branch_masks_1[soc1.core.rob.io_commit_uops_0_rob_idx] == 12'b0 : 1'b1) &&
	  (soc1.core.rob.will_commit_1 ? (rob_branch_masks_1[{soc1.core.rob.rob_head, 1'b1}] == 12'b0) && rob_branch_masks_1[soc1.core.rob.io_commit_uops_1_rob_idx] == 12'b0 : 1'b1)
	;

	//function that returns true if the given ID in store queue is above or equal stq_head and below stq_tail
	function automatic isInBoundsSTQ_1;
	//4-bit ID of the store queue entry
	input [3:0] id;
	begin
	//distinguish between positions of head and tail
	if (soc1.lsu.stq_head < soc1.lsu.stq_tail)
	begin
	  isInBoundsSTQ_1 =  id >= soc1.lsu.stq_head && id < soc1.lsu.stq_tail;
	end
	else if (soc1.lsu.stq_head > soc1.lsu.stq_tail)
	begin
	  isInBoundsSTQ_1 = id >= soc1.lsu.stq_head || id < soc1.lsu.stq_tail;
	end
	else // soc1.lsu.stq_head == soc1.lsu.stq_tail
	begin
	  isInBoundsSTQ_1 = 1'b1; // stq is full or empty, handled separately
	end
	end
	endfunction

	//stores that are not inside FIFO bounds have to be invalid to avoid unreachable dependencies
	wire stq_check_invalidated_entries_1;
	assign stq_check_invalidated_entries_1 =
	//check if misprediction happened last cycle
	  (soc1.core.b2_mispredict
	    ?
	    (isInBoundsSTQ_1(4'h0) && ROBisOlder(soc1.lsu.stq_0_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_0_valid : !soc1.lsu.stq_0_valid || soc1.lsu.stq_0_bits_committed) &&
	    (isInBoundsSTQ_1(4'h1) && ROBisOlder(soc1.lsu.stq_1_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_1_valid : !soc1.lsu.stq_1_valid || soc1.lsu.stq_1_bits_committed) &&
	    (isInBoundsSTQ_1(4'h2) && ROBisOlder(soc1.lsu.stq_2_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_2_valid : !soc1.lsu.stq_2_valid || soc1.lsu.stq_2_bits_committed) &&
	    (isInBoundsSTQ_1(4'h3) && ROBisOlder(soc1.lsu.stq_3_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_3_valid : !soc1.lsu.stq_3_valid || soc1.lsu.stq_3_bits_committed) &&
	    (isInBoundsSTQ_1(4'h4) && ROBisOlder(soc1.lsu.stq_4_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_4_valid : !soc1.lsu.stq_4_valid || soc1.lsu.stq_4_bits_committed) &&
	    (isInBoundsSTQ_1(4'h5) && ROBisOlder(soc1.lsu.stq_5_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_5_valid : !soc1.lsu.stq_5_valid || soc1.lsu.stq_5_bits_committed) &&
	    (isInBoundsSTQ_1(4'h6) && ROBisOlder(soc1.lsu.stq_6_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_6_valid : !soc1.lsu.stq_6_valid || soc1.lsu.stq_6_bits_committed) &&
	    (isInBoundsSTQ_1(4'h7) && ROBisOlder(soc1.lsu.stq_7_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_7_valid : !soc1.lsu.stq_7_valid || soc1.lsu.stq_7_bits_committed) &&
	    (isInBoundsSTQ_1(4'h8) && ROBisOlder(soc1.lsu.stq_8_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_8_valid : !soc1.lsu.stq_8_valid || soc1.lsu.stq_8_bits_committed) &&
	    (isInBoundsSTQ_1(4'h9) && ROBisOlder(soc1.lsu.stq_9_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_9_valid : !soc1.lsu.stq_9_valid || soc1.lsu.stq_9_bits_committed) &&
	    (isInBoundsSTQ_1(4'ha) && ROBisOlder(soc1.lsu.stq_10_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_10_valid : !soc1.lsu.stq_10_valid || soc1.lsu.stq_10_bits_committed) &&
	    (isInBoundsSTQ_1(4'hb) && ROBisOlder(soc1.lsu.stq_11_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_11_valid : !soc1.lsu.stq_11_valid || soc1.lsu.stq_11_bits_committed) &&
	    (isInBoundsSTQ_1(4'hc) && ROBisOlder(soc1.lsu.stq_12_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_12_valid : !soc1.lsu.stq_12_valid || soc1.lsu.stq_12_bits_committed) &&
	    (isInBoundsSTQ_1(4'hd) && ROBisOlder(soc1.lsu.stq_13_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_13_valid : !soc1.lsu.stq_13_valid || soc1.lsu.stq_13_bits_committed) &&
	    (isInBoundsSTQ_1(4'he) && ROBisOlder(soc1.lsu.stq_14_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_14_valid : !soc1.lsu.stq_14_valid || soc1.lsu.stq_14_bits_committed) &&
	    (isInBoundsSTQ_1(4'hf) && ROBisOlder(soc1.lsu.stq_15_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.stq_15_valid : !soc1.lsu.stq_15_valid || soc1.lsu.stq_15_bits_committed)
	    :
				//check if stq is empty, full or none of both
				((soc1.lsu.stq_head == soc1.lsu.stq_tail)
				?
					(soc1.lsu.stq_0_valid | soc1.lsu.stq_1_valid | soc1.lsu.stq_2_valid | soc1.lsu.stq_3_valid | soc1.lsu.stq_4_valid | soc1.lsu.stq_5_valid |	soc1.lsu.stq_6_valid | soc1.lsu.stq_7_valid | soc1.lsu.stq_8_valid | soc1.lsu.stq_12_valid | soc1.lsu.stq_13_valid | soc1.lsu.stq_14_valid | soc1.lsu.stq_15_valid)
					 == 1'b1
					 ?
				 		//if one is valid, stq has to be full
						(soc1.lsu.stq_0_valid & soc1.lsu.stq_1_valid & soc1.lsu.stq_2_valid &
						soc1.lsu.stq_3_valid & soc1.lsu.stq_4_valid & soc1.lsu.stq_5_valid &
						soc1.lsu.stq_6_valid & soc1.lsu.stq_7_valid & soc1.lsu.stq_8_valid &
						soc1.lsu.stq_9_valid & soc1.lsu.stq_10_valid & soc1.lsu.stq_11_valid &
						soc1.lsu.stq_12_valid & soc1.lsu.stq_13_valid & soc1.lsu.stq_14_valid &
						soc1.lsu.stq_15_valid) == 1'b1
					 :
						//if equal stq is empty
						(soc1.lsu.stq_0_valid | soc1.lsu.stq_1_valid | soc1.lsu.stq_2_valid |
						soc1.lsu.stq_3_valid | soc1.lsu.stq_4_valid | soc1.lsu.stq_5_valid |
						soc1.lsu.stq_6_valid | soc1.lsu.stq_7_valid | soc1.lsu.stq_8_valid |
						soc1.lsu.stq_9_valid | soc1.lsu.stq_10_valid | soc1.lsu.stq_11_valid |
						soc1.lsu.stq_12_valid | soc1.lsu.stq_13_valid | soc1.lsu.stq_14_valid |
						soc1.lsu.stq_15_valid) == 1'b0
				:
					//if not empty and not full, only valid bits with ID greater equal head or less than tail are set
					(isInBoundsSTQ_1(4'h0) ? soc1.lsu.stq_0_valid : !soc1.lsu.stq_0_valid) &&
					(isInBoundsSTQ_1(4'h1) ? soc1.lsu.stq_1_valid : !soc1.lsu.stq_1_valid) &&
					(isInBoundsSTQ_1(4'h2) ? soc1.lsu.stq_2_valid : !soc1.lsu.stq_2_valid) &&
					(isInBoundsSTQ_1(4'h3) ? soc1.lsu.stq_3_valid : !soc1.lsu.stq_3_valid) &&
					(isInBoundsSTQ_1(4'h4) ? soc1.lsu.stq_4_valid : !soc1.lsu.stq_4_valid) &&
					(isInBoundsSTQ_1(4'h5) ? soc1.lsu.stq_5_valid : !soc1.lsu.stq_5_valid) &&
					(isInBoundsSTQ_1(4'h6) ? soc1.lsu.stq_6_valid : !soc1.lsu.stq_6_valid) &&
					(isInBoundsSTQ_1(4'h7) ? soc1.lsu.stq_7_valid : !soc1.lsu.stq_7_valid) &&
					(isInBoundsSTQ_1(4'h8) ? soc1.lsu.stq_8_valid : !soc1.lsu.stq_8_valid) &&
					(isInBoundsSTQ_1(4'h9) ? soc1.lsu.stq_9_valid : !soc1.lsu.stq_9_valid) &&
					(isInBoundsSTQ_1(4'ha) ? soc1.lsu.stq_10_valid : !soc1.lsu.stq_10_valid) &&
					(isInBoundsSTQ_1(4'hb) ? soc1.lsu.stq_11_valid : !soc1.lsu.stq_11_valid) &&
					(isInBoundsSTQ_1(4'hc) ? soc1.lsu.stq_12_valid : !soc1.lsu.stq_12_valid) &&
					(isInBoundsSTQ_1(4'hd) ? soc1.lsu.stq_13_valid : !soc1.lsu.stq_13_valid) &&
					(isInBoundsSTQ_1(4'he) ? soc1.lsu.stq_14_valid : !soc1.lsu.stq_14_valid) &&
					(isInBoundsSTQ_1(4'hf) ? soc1.lsu.stq_15_valid : !soc1.lsu.stq_15_valid)
	  			)
	);

	//function that returns true if the given ID in load queue is above or equal ldq_head and below ldq_tail
	function automatic isInBoundsLDQ_1;
	  //4-bit ID of the load queue entry
	  input [3:0] id;
	  begin
	    //distinguish between positions of head and tail
	    if (soc1.lsu.ldq_head < soc1.lsu.ldq_tail)
	    begin
	      isInBoundsLDQ_1 =  id >= soc1.lsu.ldq_head && id < soc1.lsu.ldq_tail;
	    end
	    else if (soc1.lsu.ldq_head > soc1.lsu.ldq_tail)
	    begin
	      isInBoundsLDQ_1 = id >= soc1.lsu.ldq_head || id < soc1.lsu.ldq_tail;
	    end
	    else // soc1.lsu.ldq_head == soc1.lsu.ldq_tail
	    begin
	      isInBoundsLDQ_1 = 1'b1; // ldq is full or empty, handled separately
	    end
	  end
	endfunction

	//loads that are not inside FIFO bounds have to be invalid to avoid unreachable dependencies
	wire ldq_check_invalidated_entries_1;
	assign ldq_check_invalidated_entries_1 =
	//check if misprediction happened last cycle
		soc1.core.b2_mispredict
		?
			(isInBoundsLDQ_1(4'h0) && ROBisOlder(soc1.lsu.ldq_0_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_0_valid : !soc1.lsu.ldq_0_valid) &&
			(isInBoundsLDQ_1(4'h1) && ROBisOlder(soc1.lsu.ldq_1_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_1_valid : !soc1.lsu.ldq_1_valid) &&
			(isInBoundsLDQ_1(4'h2) && ROBisOlder(soc1.lsu.ldq_2_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_2_valid : !soc1.lsu.ldq_2_valid) &&
			(isInBoundsLDQ_1(4'h3) && ROBisOlder(soc1.lsu.ldq_3_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_3_valid : !soc1.lsu.ldq_3_valid) &&
			(isInBoundsLDQ_1(4'h4) && ROBisOlder(soc1.lsu.ldq_4_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_4_valid : !soc1.lsu.ldq_4_valid) &&
			(isInBoundsLDQ_1(4'h5) && ROBisOlder(soc1.lsu.ldq_5_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_5_valid : !soc1.lsu.ldq_5_valid) &&
			(isInBoundsLDQ_1(4'h6) && ROBisOlder(soc1.lsu.ldq_6_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_6_valid : !soc1.lsu.ldq_6_valid) &&
			(isInBoundsLDQ_1(4'h7) && ROBisOlder(soc1.lsu.ldq_7_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_7_valid : !soc1.lsu.ldq_7_valid) &&
			(isInBoundsLDQ_1(4'h8) && ROBisOlder(soc1.lsu.ldq_8_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_8_valid : !soc1.lsu.ldq_8_valid) &&
			(isInBoundsLDQ_1(4'h9) && ROBisOlder(soc1.lsu.ldq_9_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_9_valid : !soc1.lsu.ldq_9_valid) &&
			(isInBoundsLDQ_1(4'ha) && ROBisOlder(soc1.lsu.ldq_10_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_10_valid : !soc1.lsu.ldq_10_valid) &&
			(isInBoundsLDQ_1(4'hb) && ROBisOlder(soc1.lsu.ldq_11_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_11_valid : !soc1.lsu.ldq_11_valid) &&
			(isInBoundsLDQ_1(4'hc) && ROBisOlder(soc1.lsu.ldq_12_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_12_valid : !soc1.lsu.ldq_12_valid) &&
			(isInBoundsLDQ_1(4'hd) && ROBisOlder(soc1.lsu.ldq_13_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_13_valid : !soc1.lsu.ldq_13_valid) &&
			(isInBoundsLDQ_1(4'he) && ROBisOlder(soc1.lsu.ldq_14_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_14_valid : !soc1.lsu.ldq_14_valid) &&
			(isInBoundsLDQ_1(4'hf) && ROBisOlder(soc1.lsu.ldq_15_bits_uop_rob_idx, soc1.core.b2_uop_rob_idx, soc1.core.rob.io_rob_head_idx) ? soc1.lsu.ldq_15_valid : !soc1.lsu.ldq_15_valid)
		:
			//if equal ldq is empty
			(soc1.lsu.ldq_head == soc1.lsu.ldq_tail
			?
		 		(soc1.lsu.ldq_0_valid | soc1.lsu.ldq_1_valid | soc1.lsu.ldq_2_valid | soc1.lsu.ldq_3_valid | soc1.lsu.ldq_4_valid | soc1.lsu.ldq_5_valid |	soc1.lsu.ldq_6_valid | soc1.lsu.ldq_7_valid | soc1.lsu.ldq_8_valid | soc1.lsu.ldq_12_valid | soc1.lsu.ldq_13_valid | soc1.lsu.ldq_14_valid | soc1.lsu.ldq_15_valid)
				 == 1'b1
				?
					//if one is valid, ldq has to be full
					(soc1.lsu.ldq_0_valid & soc1.lsu.ldq_1_valid & soc1.lsu.ldq_2_valid &
					soc1.lsu.ldq_3_valid & soc1.lsu.ldq_4_valid & soc1.lsu.ldq_5_valid &
					soc1.lsu.ldq_6_valid & soc1.lsu.ldq_7_valid & soc1.lsu.ldq_8_valid &
					soc1.lsu.ldq_9_valid & soc1.lsu.ldq_10_valid & soc1.lsu.ldq_11_valid &
					soc1.lsu.ldq_12_valid & soc1.lsu.ldq_13_valid & soc1.lsu.ldq_14_valid &
					soc1.lsu.ldq_15_valid) == 1'b1
				:
					//if empty all valid bits are zero
					(soc1.lsu.ldq_0_valid | soc1.lsu.ldq_1_valid | soc1.lsu.ldq_2_valid |
					soc1.lsu.ldq_3_valid | soc1.lsu.ldq_4_valid | soc1.lsu.ldq_5_valid |
					soc1.lsu.ldq_6_valid | soc1.lsu.ldq_7_valid | soc1.lsu.ldq_8_valid |
					soc1.lsu.ldq_9_valid | soc1.lsu.ldq_10_valid | soc1.lsu.ldq_11_valid |
					soc1.lsu.ldq_12_valid | soc1.lsu.ldq_13_valid | soc1.lsu.ldq_14_valid |
					soc1.lsu.ldq_15_valid) == 1'b0
			:
				//if not empty and not full, only valid bits with ID greater equal head or less than tail are set
				(isInBoundsLDQ_1(4'h0) ? soc1.lsu.ldq_0_valid : !soc1.lsu.ldq_0_valid) &&
				(isInBoundsLDQ_1(4'h1) ? soc1.lsu.ldq_1_valid : !soc1.lsu.ldq_1_valid) &&
				(isInBoundsLDQ_1(4'h2) ? soc1.lsu.ldq_2_valid : !soc1.lsu.ldq_2_valid) &&
				(isInBoundsLDQ_1(4'h3) ? soc1.lsu.ldq_3_valid : !soc1.lsu.ldq_3_valid) &&
				(isInBoundsLDQ_1(4'h4) ? soc1.lsu.ldq_4_valid : !soc1.lsu.ldq_4_valid) &&
				(isInBoundsLDQ_1(4'h5) ? soc1.lsu.ldq_5_valid : !soc1.lsu.ldq_5_valid) &&
				(isInBoundsLDQ_1(4'h6) ? soc1.lsu.ldq_6_valid : !soc1.lsu.ldq_6_valid) &&
				(isInBoundsLDQ_1(4'h7) ? soc1.lsu.ldq_7_valid : !soc1.lsu.ldq_7_valid) &&
				(isInBoundsLDQ_1(4'h8) ? soc1.lsu.ldq_8_valid : !soc1.lsu.ldq_8_valid) &&
				(isInBoundsLDQ_1(4'h9) ? soc1.lsu.ldq_9_valid : !soc1.lsu.ldq_9_valid) &&
				(isInBoundsLDQ_1(4'ha) ? soc1.lsu.ldq_10_valid : !soc1.lsu.ldq_10_valid) &&
				(isInBoundsLDQ_1(4'hb) ? soc1.lsu.ldq_11_valid : !soc1.lsu.ldq_11_valid) &&
				(isInBoundsLDQ_1(4'hc) ? soc1.lsu.ldq_12_valid : !soc1.lsu.ldq_12_valid) &&
				(isInBoundsLDQ_1(4'hd) ? soc1.lsu.ldq_13_valid : !soc1.lsu.ldq_13_valid) &&
				(isInBoundsLDQ_1(4'he) ? soc1.lsu.ldq_14_valid : !soc1.lsu.ldq_14_valid) &&
				(isInBoundsLDQ_1(4'hf) ? soc1.lsu.ldq_15_valid : !soc1.lsu.ldq_15_valid)
			)
	;

	wire consistent_buffer_br_masks_1;
	assign consistent_buffer_br_masks_1 =
	  (soc1.core.csr_exe_unit.alu.r_valids_0 ? rob_valids_1[soc1.core.csr_exe_unit.alu.r_uops_0_rob_idx] && soc1.core.csr_exe_unit.alu.r_uops_0_br_mask == rob_branch_masks_1[soc1.core.csr_exe_unit.alu.r_uops_0_rob_idx] : 1'b1) &&
	  ((soc1.core.csr_exe_unit.div.div.state == 3'h3) ||(soc1.core.csr_exe_unit.div.div.state == 3'h7) ? rob_valids_1[soc1.core.csr_exe_unit.div.r_uop_rob_idx] && soc1.core.csr_exe_unit.div.r_uop_br_mask == rob_branch_masks_1[soc1.core.csr_exe_unit.div.r_uop_rob_idx] : 1'b1) &&
	  (soc1.core.iregister_read.exe_reg_valids_0  /*&& !(soc1.core.iregister_read.exe_reg_uops_0_uses_stq && stq_committed_1[soc1.core.iregister_read.exe_reg_uops_0_stq_idx]) */? rob_valids_1[soc1.core.iregister_read.exe_reg_uops_0_rob_idx] && soc1.core.iregister_read.exe_reg_uops_0_br_mask == rob_branch_masks_1[soc1.core.iregister_read.exe_reg_uops_0_rob_idx] : 1'b1) &&
	  (soc1.core.iregister_read.exe_reg_valids_1  /*&& !(soc1.core.iregister_read.exe_reg_uops_1_uses_stq && stq_committed_1[soc1.core.iregister_read.exe_reg_uops_1_stq_idx]) */? rob_valids_1[soc1.core.iregister_read.exe_reg_uops_1_rob_idx] && soc1.core.iregister_read.exe_reg_uops_1_br_mask == rob_branch_masks_1[soc1.core.iregister_read.exe_reg_uops_1_rob_idx] : 1'b1) &&
	  (soc1.core.iregister_read.exe_reg_valids_2  /*&& !(soc1.core.iregister_read.exe_reg_uops_2_uses_stq && stq_committed_1[soc1.core.iregister_read.exe_reg_uops_2_stq_idx]) */? rob_valids_1[soc1.core.iregister_read.exe_reg_uops_2_rob_idx] && soc1.core.iregister_read.exe_reg_uops_2_br_mask == rob_branch_masks_1[soc1.core.iregister_read.exe_reg_uops_2_rob_idx] : 1'b1) &&
	  (soc1.core.iregister_read.rrd_valids_0_REG  /*&& !(soc1.core.iregister_read.rrd_uops_0_REG_uses_stq && stq_committed_1[soc1.core.iregister_read.rrd_uops_0_REG_stq_idx]) */? rob_valids_1[soc1.core.iregister_read.rrd_uops_0_REG_rob_idx] && soc1.core.iregister_read.rrd_uops_0_REG_br_mask == rob_branch_masks_1[soc1.core.iregister_read.rrd_uops_0_REG_rob_idx] : 1'b1) &&
	  (soc1.core.iregister_read.rrd_valids_1_REG  /*&& !(soc1.core.iregister_read.rrd_uops_1_REG_uses_stq && stq_committed_1[soc1.core.iregister_read.rrd_uops_1_REG_stq_idx]) */? rob_valids_1[soc1.core.iregister_read.rrd_uops_1_REG_rob_idx] && soc1.core.iregister_read.rrd_uops_1_REG_br_mask == rob_branch_masks_1[soc1.core.iregister_read.rrd_uops_1_REG_rob_idx] : 1'b1) &&
	  (soc1.core.iregister_read.rrd_valids_2_REG  /*&& !(soc1.core.iregister_read.rrd_uops_2_REG_uses_stq && stq_committed_1[soc1.core.iregister_read.rrd_uops_2_REG_stq_idx]) */? rob_valids_1[soc1.core.iregister_read.rrd_uops_2_REG_rob_idx] && soc1.core.iregister_read.rrd_uops_2_REG_br_mask == rob_branch_masks_1[soc1.core.iregister_read.rrd_uops_2_REG_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.queue.valids_0 ? rob_valids_1[soc1.core.jmp_unit.queue.uops_0_rob_idx] && soc1.core.jmp_unit.queue.uops_0_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.queue.uops_0_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.queue.valids_1 ? rob_valids_1[soc1.core.jmp_unit.queue.uops_1_rob_idx] && soc1.core.jmp_unit.queue.uops_1_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.queue.uops_1_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.queue.valids_2 ? rob_valids_1[soc1.core.jmp_unit.queue.uops_2_rob_idx] && soc1.core.jmp_unit.queue.uops_2_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.queue.uops_2_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.queue.valids_3 ? rob_valids_1[soc1.core.jmp_unit.queue.uops_3_rob_idx] && soc1.core.jmp_unit.queue.uops_3_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.queue.uops_3_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.queue.valids_4 ? rob_valids_1[soc1.core.jmp_unit.queue.uops_4_rob_idx] && soc1.core.jmp_unit.queue.uops_4_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.queue.uops_4_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.alu.r_valids_0 ? rob_valids_1[soc1.core.jmp_unit.alu.r_uops_0_rob_idx] && soc1.core.jmp_unit.alu.r_uops_0_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.alu.r_uops_0_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.alu.r_valids_1 ? rob_valids_1[soc1.core.jmp_unit.alu.r_uops_1_rob_idx] && soc1.core.jmp_unit.alu.r_uops_1_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.alu.r_uops_1_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.alu.r_valids_2 ? rob_valids_1[soc1.core.jmp_unit.alu.r_uops_2_rob_idx] && soc1.core.jmp_unit.alu.r_uops_2_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.alu.r_uops_2_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.ifpu.r_valids_0 ? rob_valids_1[soc1.core.jmp_unit.ifpu.r_uops_0_rob_idx] && soc1.core.jmp_unit.ifpu.r_uops_0_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.ifpu.r_uops_0_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.ifpu.r_valids_1 ? rob_valids_1[soc1.core.jmp_unit.ifpu.r_uops_1_rob_idx] && soc1.core.jmp_unit.ifpu.r_uops_1_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.ifpu.r_uops_1_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.imul.r_valids_0 ? rob_valids_1[soc1.core.jmp_unit.imul.r_uops_0_rob_idx] && soc1.core.jmp_unit.imul.r_uops_0_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.imul.r_uops_0_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.imul.r_valids_1 ? rob_valids_1[soc1.core.jmp_unit.imul.r_uops_1_rob_idx] && soc1.core.jmp_unit.imul.r_uops_1_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.imul.r_uops_1_rob_idx] : 1'b1) &&
	  (soc1.core.jmp_unit.imul.r_valids_2 ? rob_valids_1[soc1.core.jmp_unit.imul.r_uops_2_rob_idx] && soc1.core.jmp_unit.imul.r_uops_2_br_mask == rob_branch_masks_1[soc1.core.jmp_unit.imul.r_uops_2_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_0.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_1.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_2.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_3.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_4.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_5.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_6.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_7.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_8.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_9.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_10.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_11.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_12.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_13.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_14.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fp_issue_unit.slots_15.io_valid /*&& !(soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx] && soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.queue.valids_0 /*&& !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.queue.valids_1 /*&& !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.queue.valids_2 /*&& !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.queue.valids_3 /*&& !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.queue.valids_4 /*&& !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.queue.valids_5 /*&& !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.queue.valids_6 /*&& !(soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0 ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1 ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2 ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_val ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_val ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_0 && !(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_stq_idx]) ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_1 && !(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_stq_idx]) ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_2 && !(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_stq_idx]) ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_3 && !(soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_stq_idx]) ? rob_valids_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx] && soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fregister_read.exe_reg_valids_0 /*&& !(soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx] && soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx] : 1'b1) &&
	  (soc1.core.fp_pipeline.fregister_read.rrd_valids_0_REG /*&& !(soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_stq_idx]) */? rob_valids_1[soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx] && soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_br_mask == rob_branch_masks_1[soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_0.io_valid /*&& !(soc1.core.int_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_0.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_0.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_0.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_0.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_1.io_valid /*&& !(soc1.core.int_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_1.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_1.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_1.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_1.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_2.io_valid /*&& !(soc1.core.int_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_2.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_2.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_2.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_2.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_3.io_valid /*&& !(soc1.core.int_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_3.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_3.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_3.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_3.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_4.io_valid /*&& !(soc1.core.int_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_4.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_4.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_4.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_4.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_5.io_valid /*&& !(soc1.core.int_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_5.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_5.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_5.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_5.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_6.io_valid /*&& !(soc1.core.int_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_6.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_6.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_6.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_6.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_7.io_valid /*&& !(soc1.core.int_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_7.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_7.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_7.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_7.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_8.io_valid /*&& !(soc1.core.int_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_8.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_8.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_8.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_8.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_9.io_valid /*&& !(soc1.core.int_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_9.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_9.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_9.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_9.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_10.io_valid /*&& !(soc1.core.int_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_10.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_10.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_10.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_10.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_11.io_valid /*&& !(soc1.core.int_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_11.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_11.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_11.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_11.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_12.io_valid /*&& !(soc1.core.int_issue_unit.slots_12.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_12.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_12.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_12.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_12.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_13.io_valid /*&& !(soc1.core.int_issue_unit.slots_13.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_13.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_13.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_13.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_13.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_14.io_valid /*&& !(soc1.core.int_issue_unit.slots_14.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_14.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_14.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_14.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_14.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_15.io_valid /*&& !(soc1.core.int_issue_unit.slots_15.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_15.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_15.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_15.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_15.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_16.io_valid /*&& !(soc1.core.int_issue_unit.slots_16.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_16.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_16.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_16.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_16.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_17.io_valid /*&& !(soc1.core.int_issue_unit.slots_17.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_17.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_17.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_17.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_17.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_18.io_valid /*&& !(soc1.core.int_issue_unit.slots_18.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_18.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_18.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_18.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_18.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.int_issue_unit.slots_19.io_valid /*&& !(soc1.core.int_issue_unit.slots_19.slot_uop_uses_stq && stq_committed_1[soc1.core.int_issue_unit.slots_19.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.int_issue_unit.slots_19.slot_uop_rob_idx] && soc1.core.int_issue_unit.slots_19.slot_uop_br_mask == rob_branch_masks_1[soc1.core.int_issue_unit.slots_19.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_0.io_valid /*&& !(soc1.core.mem_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_0.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_0.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_0.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_0.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_1.io_valid /*&& !(soc1.core.mem_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_1.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_1.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_1.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_1.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_2.io_valid /*&& !(soc1.core.mem_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_2.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_2.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_2.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_2.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_3.io_valid /*&& !(soc1.core.mem_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_3.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_3.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_3.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_3.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_4.io_valid /*&& !(soc1.core.mem_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_4.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_4.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_4.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_4.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_5.io_valid /*&& !(soc1.core.mem_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_5.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_5.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_5.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_5.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_6.io_valid /*&& !(soc1.core.mem_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_6.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_6.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_6.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_6.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_7.io_valid /*&& !(soc1.core.mem_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_7.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_7.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_7.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_7.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_8.io_valid /*&& !(soc1.core.mem_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_8.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_8.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_8.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_8.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_9.io_valid /*&& !(soc1.core.mem_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_9.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_9.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_9.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_9.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_10.io_valid /*&& !(soc1.core.mem_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_10.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_10.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_10.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_10.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.core.mem_issue_unit.slots_11.io_valid /*&& !(soc1.core.mem_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_1[soc1.core.mem_issue_unit.slots_11.slot_uop_stq_idx]) */? rob_valids_1[soc1.core.mem_issue_unit.slots_11.slot_uop_rob_idx] && soc1.core.mem_issue_unit.slots_11.slot_uop_br_mask == rob_branch_masks_1[soc1.core.mem_issue_unit.slots_11.slot_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_0_valid ? rob_valids_1[soc1.lsu.ldq_0_bits_uop_rob_idx] && soc1.lsu.ldq_0_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_0_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_1_valid ? rob_valids_1[soc1.lsu.ldq_1_bits_uop_rob_idx] && soc1.lsu.ldq_1_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_1_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_2_valid ? rob_valids_1[soc1.lsu.ldq_2_bits_uop_rob_idx] && soc1.lsu.ldq_2_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_2_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_3_valid ? rob_valids_1[soc1.lsu.ldq_3_bits_uop_rob_idx] && soc1.lsu.ldq_3_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_3_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_4_valid ? rob_valids_1[soc1.lsu.ldq_4_bits_uop_rob_idx] && soc1.lsu.ldq_4_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_4_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_5_valid ? rob_valids_1[soc1.lsu.ldq_5_bits_uop_rob_idx] && soc1.lsu.ldq_5_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_5_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_6_valid ? rob_valids_1[soc1.lsu.ldq_6_bits_uop_rob_idx] && soc1.lsu.ldq_6_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_6_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_7_valid ? rob_valids_1[soc1.lsu.ldq_7_bits_uop_rob_idx] && soc1.lsu.ldq_7_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_7_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_8_valid ? rob_valids_1[soc1.lsu.ldq_8_bits_uop_rob_idx] && soc1.lsu.ldq_8_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_8_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_9_valid ? rob_valids_1[soc1.lsu.ldq_9_bits_uop_rob_idx] && soc1.lsu.ldq_9_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_9_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_10_valid ? rob_valids_1[soc1.lsu.ldq_10_bits_uop_rob_idx] && soc1.lsu.ldq_10_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_10_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_11_valid ? rob_valids_1[soc1.lsu.ldq_11_bits_uop_rob_idx] && soc1.lsu.ldq_11_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_11_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_12_valid ? rob_valids_1[soc1.lsu.ldq_12_bits_uop_rob_idx] && soc1.lsu.ldq_12_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_12_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_13_valid ? rob_valids_1[soc1.lsu.ldq_13_bits_uop_rob_idx] && soc1.lsu.ldq_13_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_13_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_14_valid ? rob_valids_1[soc1.lsu.ldq_14_bits_uop_rob_idx] && soc1.lsu.ldq_14_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_14_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_15_valid ? rob_valids_1[soc1.lsu.ldq_15_bits_uop_rob_idx] && soc1.lsu.ldq_15_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.ldq_15_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.fired_sfence_0 ? rob_valids_1[soc1.lsu.mem_incoming_uop_0_rob_idx] && soc1.lsu.mem_incoming_uop_0_br_mask == rob_branch_masks_1[soc1.lsu.mem_incoming_uop_0_rob_idx] : 1'b1) &&
	  ((soc1.lsu.fired_stad_incoming_REG || soc1.lsu.fired_sta_incoming_REG || soc1.lsu.fired_std_incoming_REG) /*&& !stq_committed_1[soc1.lsu.mem_stq_incoming_e_0_bits_uop_stq_idx] */? rob_valids_1[soc1.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx] && soc1.lsu.mem_stq_incoming_e_0_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.fired_sta_retry_REG /*&& !stq_committed_1[soc1.lsu.mem_stq_retry_e_bits_uop_stq_idx] */? rob_valids_1[soc1.lsu.mem_stq_retry_e_bits_uop_rob_idx] && soc1.lsu.mem_stq_retry_e_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.mem_stq_retry_e_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.mem_xcpt_valids_0 /*&& !(soc1.lsu.mem_xcpt_uops_0_uses_stq && stq_committed_1[soc1.lsu.mem_xcpt_uops_0_stq_idx]) */? rob_valids_1[soc1.lsu.mem_xcpt_uops_0_rob_idx] && soc1.lsu.mem_xcpt_uops_0_br_mask == rob_branch_masks_1[soc1.lsu.mem_xcpt_uops_0_rob_idx] : 1'b1) &&
	  (soc1.lsu.fired_stdf_incoming /*&& !stq_committed_1[soc1.lsu.mem_stdf_uop_stq_idx] */? rob_valids_1[soc1.lsu.mem_stdf_uop_rob_idx] && soc1.lsu.mem_stdf_uop_br_mask == rob_branch_masks_1[soc1.lsu.mem_stdf_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stdf_clr_bsy_valid ? rob_valids_1[soc1.lsu.stdf_clr_bsy_rob_idx] && soc1.lsu.stdf_clr_bsy_brmask == rob_branch_masks_1[soc1.lsu.stdf_clr_bsy_rob_idx] : 1'b1) &&
	  //stores do not have to be checked after they are committed (their ROB entry can be used for another uop then)
	  (soc1.lsu.stq_0_valid && !soc1.lsu.stq_0_bits_committed ? rob_valids_1[soc1.lsu.stq_0_bits_uop_rob_idx] && soc1.lsu.stq_0_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_0_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_1_valid && !soc1.lsu.stq_1_bits_committed ? rob_valids_1[soc1.lsu.stq_1_bits_uop_rob_idx] && soc1.lsu.stq_1_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_1_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_2_valid && !soc1.lsu.stq_2_bits_committed ? rob_valids_1[soc1.lsu.stq_2_bits_uop_rob_idx] && soc1.lsu.stq_2_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_2_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_3_valid && !soc1.lsu.stq_3_bits_committed ? rob_valids_1[soc1.lsu.stq_3_bits_uop_rob_idx] && soc1.lsu.stq_3_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_3_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_4_valid && !soc1.lsu.stq_4_bits_committed ? rob_valids_1[soc1.lsu.stq_4_bits_uop_rob_idx] && soc1.lsu.stq_4_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_4_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_5_valid && !soc1.lsu.stq_5_bits_committed ? rob_valids_1[soc1.lsu.stq_5_bits_uop_rob_idx] && soc1.lsu.stq_5_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_5_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_6_valid && !soc1.lsu.stq_6_bits_committed ? rob_valids_1[soc1.lsu.stq_6_bits_uop_rob_idx] && soc1.lsu.stq_6_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_6_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_7_valid && !soc1.lsu.stq_7_bits_committed ? rob_valids_1[soc1.lsu.stq_7_bits_uop_rob_idx] && soc1.lsu.stq_7_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_7_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_8_valid && !soc1.lsu.stq_8_bits_committed ? rob_valids_1[soc1.lsu.stq_8_bits_uop_rob_idx] && soc1.lsu.stq_8_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_8_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_9_valid && !soc1.lsu.stq_9_bits_committed ? rob_valids_1[soc1.lsu.stq_9_bits_uop_rob_idx] && soc1.lsu.stq_9_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_9_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_10_valid && !soc1.lsu.stq_10_bits_committed ? rob_valids_1[soc1.lsu.stq_10_bits_uop_rob_idx] && soc1.lsu.stq_10_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_10_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_11_valid && !soc1.lsu.stq_11_bits_committed ? rob_valids_1[soc1.lsu.stq_11_bits_uop_rob_idx] && soc1.lsu.stq_11_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_11_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_12_valid && !soc1.lsu.stq_12_bits_committed ? rob_valids_1[soc1.lsu.stq_12_bits_uop_rob_idx] && soc1.lsu.stq_12_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_12_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_13_valid && !soc1.lsu.stq_13_bits_committed ? rob_valids_1[soc1.lsu.stq_13_bits_uop_rob_idx] && soc1.lsu.stq_13_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_13_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_14_valid && !soc1.lsu.stq_14_bits_committed ? rob_valids_1[soc1.lsu.stq_14_bits_uop_rob_idx] && soc1.lsu.stq_14_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_14_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.stq_15_valid && !soc1.lsu.stq_15_bits_committed ? rob_valids_1[soc1.lsu.stq_15_bits_uop_rob_idx] && soc1.lsu.stq_15_bits_uop_br_mask == rob_branch_masks_1[soc1.lsu.stq_15_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.clr_bsy_valid_0 ? rob_valids_1[soc1.lsu.clr_bsy_rob_idx_0] && soc1.lsu.clr_bsy_brmask_0 == rob_branch_masks_1[soc1.lsu.clr_bsy_rob_idx_0] : 1'b1) &&
	  (soc1.lsu.r_xcpt_valid ? rob_valids_1[soc1.lsu.r_xcpt_uop_rob_idx] && soc1.lsu.r_xcpt_uop_br_mask == rob_branch_masks_1[soc1.lsu.r_xcpt_uop_rob_idx] : 1'b1) &&

	  (soc1.dcache.mshrs.respq.valids_0
	  ? (
	    (soc1.dcache.mshrs.respq.uops_0_uses_ldq ? rob_valids_1[ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_0_ldq_idx]] && soc1.dcache.mshrs.respq.uops_0_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_0_ldq_idx]] : 1'b1) &&
	    (soc1.dcache.mshrs.respq.uops_0_uses_stq && !stq_committed_1[soc1.dcache.mshrs.respq.uops_0_stq_idx] ? rob_valids_1[stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_0_stq_idx]] && soc1.dcache.mshrs.respq.uops_0_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_0_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.respq.valids_1
	  ? (
	    (soc1.dcache.mshrs.respq.uops_1_uses_ldq ? rob_valids_1[ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_1_ldq_idx]] && soc1.dcache.mshrs.respq.uops_1_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_1_ldq_idx]] : 1'b1) &&
	    (soc1.dcache.mshrs.respq.uops_1_uses_stq && !stq_committed_1[soc1.dcache.mshrs.respq.uops_1_stq_idx] ? rob_valids_1[stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_1_stq_idx]] && soc1.dcache.mshrs.respq.uops_1_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_1_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.respq.valids_2
	  ? (
	    (soc1.dcache.mshrs.respq.uops_2_uses_ldq ? rob_valids_1[ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_2_ldq_idx]] && soc1.dcache.mshrs.respq.uops_2_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_2_ldq_idx]] : 1'b1) &&
	    (soc1.dcache.mshrs.respq.uops_2_uses_stq && !stq_committed_1[soc1.dcache.mshrs.respq.uops_2_stq_idx] ? rob_valids_1[stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_2_stq_idx]] && soc1.dcache.mshrs.respq.uops_2_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_2_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.respq.valids_3
	  ? (
	    (soc1.dcache.mshrs.respq.uops_3_uses_ldq ? rob_valids_1[ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_3_ldq_idx]] && soc1.dcache.mshrs.respq.uops_3_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.respq.uops_3_ldq_idx]] : 1'b1) &&
	    (soc1.dcache.mshrs.respq.uops_3_uses_stq && !stq_committed_1[soc1.dcache.mshrs.respq.uops_3_stq_idx] ? rob_valids_1[stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_3_stq_idx]] && soc1.dcache.mshrs.respq.uops_3_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.respq.uops_3_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mmios_0.state != 2'b0
	  ? (
	    (soc1.dcache.mshrs.mmios_0.req_uop_uses_ldq ? rob_valids_1[ldq_rob_idx_1[soc1.dcache.mshrs.mmios_0.req_uop_ldq_idx]] && soc1.dcache.mshrs.mmios_0.req_uop_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mmios_0.req_uop_ldq_idx]] : 1'b1) &&
	    (soc1.dcache.mshrs.mmios_0.req_uop_uses_stq && !stq_committed_1[soc1.dcache.mshrs.mmios_0.req_uop_stq_idx] ? rob_valids_1[stq_rob_idx_1[soc1.dcache.mshrs.mmios_0.req_uop_stq_idx]] && soc1.dcache.mshrs.mmios_0.req_uop_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mmios_0.req_uop_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_0
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_0_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_0_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_0_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_1
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_1_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_1_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_1_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_2
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_2_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_2_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_2_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_3
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_3_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_3_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_3_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_4
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_4_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_4_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_4_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_5
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_5_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_5_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_5_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_6
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_6_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_6_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_6_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_7
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_7_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_7_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_7_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_8
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_8_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_8_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_8_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_9
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_9_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_9_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_9_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_10
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_10_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_10_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_10_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_11
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_11_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_11_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_11_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_12
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_12_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_12_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_12_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_13
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_13_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_13_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_13_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_14
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_14_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_14_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_14_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_15
	  ? (
	    (soc1.dcache.mshrs.mshrs_0.rpq.uops_15_uses_ldq ? soc1.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_15_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_0.rpq.uops_15_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx] ? soc1.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_0
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_0_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_0_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_0_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_1
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_1_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_1_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_1_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_2
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_2_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_2_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_2_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_3
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_3_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_3_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_3_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_4
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_4_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_4_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_4_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_5
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_5_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_5_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_5_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_6
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_6_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_6_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_6_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_7
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_7_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_7_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_7_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_8
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_8_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_8_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_8_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_9
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_9_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_9_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_9_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_10
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_10_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_10_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_10_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_11
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_11_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_11_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_11_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_12
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_12_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_12_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_12_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_13
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_13_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_13_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_13_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_14
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_14_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_14_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_14_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_15
	  ? (
	    (soc1.dcache.mshrs.mshrs_1.rpq.uops_15_uses_ldq ? soc1.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_15_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.mshrs.mshrs_1.rpq.uops_15_uses_stq && !stq_committed[soc1.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx] ? soc1.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.s1_valid_REG
	  ? (
	    (soc1.dcache.s1_req_0_uop_uses_ldq ? soc1.dcache.s1_req_0_uop_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.s1_req_0_uop_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.s1_req_0_uop_uses_stq ? soc1.dcache.s1_req_0_uop_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.s1_req_0_uop_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc1.dcache.s2_valid_REG
	  ? (
	    (soc1.dcache.s2_req_0_uop_uses_ldq ? soc1.dcache.s2_req_0_uop_br_mask == rob_branch_masks_1[ldq_rob_idx_1[soc1.dcache.s2_req_0_uop_ldq_idx]] : 1'b1) //&&
	    )//(soc1.dcache.s2_req_0_uop_uses_stq ? soc1.dcache.s2_req_0_uop_br_mask == rob_branch_masks_1[stq_rob_idx_1[soc1.dcache.s2_req_0_uop_stq_idx]] : 1'b1))
	  :
	    1'b1)
  	;

	//check for all issue slots:
	//if the corresponding ROB entry is invalid the state of the issue slot has to be invalid too
	wire valid_issue_slots_1;
	assign valid_issue_slots_1 =
	(!rob_valids_1[soc1.core.int_issue_unit.slots_0.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_0.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_1.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_1.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_2.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_2.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_3.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_3.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_4.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_4.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_5.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_5.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_6.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_6.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_7.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_7.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_8.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_8.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_9.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_9.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_10.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_10.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_11.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_11.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_12.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_12.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_13.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_13.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_14.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_14.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_15.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_15.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_16.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_16.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_17.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_17.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_18.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_18.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.int_issue_unit.slots_19.slot_uop_rob_idx] ? soc1.core.int_issue_unit.slots_19.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_0.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_0.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_1.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_1.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_2.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_2.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_3.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_3.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_4.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_4.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_5.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_5.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_6.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_6.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_7.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_7.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_8.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_8.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_9.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_9.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_10.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_10.state == 2'b0 : 1'b1) &&
	(!rob_valids_1[soc1.core.mem_issue_unit.slots_11.slot_uop_rob_idx] ? soc1.core.mem_issue_unit.slots_11.state == 2'b0 : 1'b1);

	//check for the branch misprediction:
	//if the prediction is valid the corresponding ROB entry must be valid too
	wire valid_mispred_idx_1;
	assign valid_mispred_idx_1 =
	(soc1.core.brinfos_0_valid ? rob_valids_1[soc1.core.brinfos_0_uop_rob_idx] : 1'b1) &&
	(soc1.core.brinfos_1_valid ? rob_valids_1[soc1.core.brinfos_1_uop_rob_idx] : 1'b1);

	//check for iregister read buffers:
	//if the buffer is valid the corresponding ROB entry must be valid too
	wire valid_iregister_read_1;
	assign valid_iregister_read_1 =
	(soc1.core.iregister_read.exe_reg_valids_1 ? rob_valids_1[soc1.core.iregister_read.exe_reg_uops_1_rob_idx] : 1'b1) &&
	(soc1.core.iregister_read.exe_reg_valids_2 ? rob_valids_1[soc1.core.iregister_read.exe_reg_uops_2_rob_idx] : 1'b1) &&
	(soc1.core.iregister_read.rrd_valids_1_REG ? rob_valids_1[soc1.core.iregister_read.rrd_uops_1_REG_rob_idx] : 1'b1) &&
	(soc1.core.iregister_read.rrd_valids_2_REG ? rob_valids_1[soc1.core.iregister_read.rrd_uops_2_REG_rob_idx] : 1'b1);

	//instruction at head must be non-speculative (br_mask == 0) if it is valid
	wire no_speculative_head_1;
	assign no_speculative_head_1 =
	  rob_valids_1[soc1.core.rob.io_rob_head_idx]? (rob_branch_masks_1[soc1.core.rob.io_rob_head_idx] == 12'b0) : 1'b1;
	  
	//ensure that valid entries are not overwritten
	wire prevent_overwriting_valid_entries_1;
	assign prevent_overwriting_valid_entries_1 = 
	  (soc1.core.rob.io_enq_valids_0 ? !rob_valids_1[{soc1.core.rob.rob_tail,1'b0}] : 1'b1) &&
	  (soc1.core.rob.io_enq_valids_1 ? !rob_valids_1[{soc1.core.rob.rob_tail,1'b1}] : 1'b1);
	  
	//ROB is never full and empty
	wire full_empty_logic_1;
	assign full_empty_logic_1 = !(soc1.core.rob.full && soc1.core.rob.empty);

	//ROB is empty equals head == tail and all valid bits are 0
	wire empty_logic_1;
	assign empty_logic_1 =
	  ((soc1.core.rob.rob_head == soc1.core.rob.rob_tail) && ((rob_valids_1[0] | rob_valids_1[1] | rob_valids_1[2] | rob_valids_1[3] | rob_valids_1[4] | rob_valids_1[5] | rob_valids_1[6] | rob_valids_1[7] | rob_valids_1[8] | rob_valids_1[9] |
	    rob_valids_1[10] | rob_valids_1[11] | rob_valids_1[12] | rob_valids_1[13] | rob_valids_1[14] | rob_valids_1[15] | rob_valids_1[16] | rob_valids_1[17] | rob_valids_1[18] | rob_valids_1[19] | 
	    rob_valids_1[20] | rob_valids_1[21] | rob_valids_1[22] | rob_valids_1[23] | rob_valids_1[24] | rob_valids_1[25] | rob_valids_1[26] | rob_valids_1[27] | rob_valids_1[28] | rob_valids_1[29] | 
	    rob_valids_1[30] | rob_valids_1[31] | rob_valids_1[32] | rob_valids_1[33] | rob_valids_1[34] | rob_valids_1[35] | rob_valids_1[36] | rob_valids_1[37] | rob_valids_1[38] | rob_valids_1[39] | 
	    rob_valids_1[40] | rob_valids_1[41] | rob_valids_1[42] | rob_valids_1[43] | rob_valids_1[44] | rob_valids_1[45] | rob_valids_1[46] | rob_valids_1[47] | rob_valids_1[48] | rob_valids_1[49] | 
	    rob_valids_1[50] | rob_valids_1[51] | rob_valids_1[52] | rob_valids_1[53] | rob_valids_1[54] | rob_valids_1[55] | rob_valids_1[56] | rob_valids_1[57] | rob_valids_1[58] | rob_valids_1[59] | 
	    rob_valids_1[60] | rob_valids_1[61] | rob_valids_1[62] | rob_valids_1[63]) == 1'b0)) == soc1.core.rob.empty;
	    
	//ROB is full equals head == tail and either one of the entrys at tail is valid or tail_lsb is not set, else rob_state is rollback
	wire full_logic_1;
	assign full_logic_1 = (soc1.core.rob.rob_head == soc1.core.rob.rob_tail && soc1.core.rob.maybe_full) == soc1.core.rob.full;
	  
	//Create array for load queue valid bits
	wire ldq_valids_1 [15:0];
	assign ldq_valids_1[0] = soc1.lsu.ldq_0_valid;
	assign ldq_valids_1[1] = soc1.lsu.ldq_1_valid;
	assign ldq_valids_1[2] = soc1.lsu.ldq_2_valid;
	assign ldq_valids_1[3] = soc1.lsu.ldq_3_valid;
	assign ldq_valids_1[4] = soc1.lsu.ldq_4_valid;
	assign ldq_valids_1[5] = soc1.lsu.ldq_5_valid;
	assign ldq_valids_1[6] = soc1.lsu.ldq_6_valid;
	assign ldq_valids_1[7] = soc1.lsu.ldq_7_valid;
	assign ldq_valids_1[8] = soc1.lsu.ldq_8_valid;
	assign ldq_valids_1[9] = soc1.lsu.ldq_9_valid;
	assign ldq_valids_1[10] = soc1.lsu.ldq_10_valid;
	assign ldq_valids_1[11] = soc1.lsu.ldq_11_valid;
	assign ldq_valids_1[12] = soc1.lsu.ldq_12_valid;
	assign ldq_valids_1[13] = soc1.lsu.ldq_13_valid;
	assign ldq_valids_1[14] = soc1.lsu.ldq_14_valid;
	assign ldq_valids_1[15] = soc1.lsu.ldq_15_valid;
	  
	wire lcam_ldq_idx_valid_1;
	assign lcam_ldq_idx_valid_1 = 
	//if a load got fired, its ldq entry has to be valid
	(soc1.lsu.fired_load_incoming_REG || soc1.lsu.fired_load_retry_REG || soc1.lsu.fired_load_wakeup_REG) && !soc1.lsu.REG_1 ? ldq_valids_1[soc1.lsu.lcam_ldq_idx_0] : 1'b1;
	
	//Create array for load queue valid bits
	wire stq_valids_1 [15:0];
	assign stq_valids_1[0] = soc1.lsu.stq_0_valid;
	assign stq_valids_1[1] = soc1.lsu.stq_1_valid;
	assign stq_valids_1[2] = soc1.lsu.stq_2_valid;
	assign stq_valids_1[3] = soc1.lsu.stq_3_valid;
	assign stq_valids_1[4] = soc1.lsu.stq_4_valid;
	assign stq_valids_1[5] = soc1.lsu.stq_5_valid;
	assign stq_valids_1[6] = soc1.lsu.stq_6_valid;
	assign stq_valids_1[7] = soc1.lsu.stq_7_valid;
	assign stq_valids_1[8] = soc1.lsu.stq_8_valid;
	assign stq_valids_1[9] = soc1.lsu.stq_9_valid;
	assign stq_valids_1[10] = soc1.lsu.stq_10_valid;
	assign stq_valids_1[11] = soc1.lsu.stq_11_valid;
	assign stq_valids_1[12] = soc1.lsu.stq_12_valid;
	assign stq_valids_1[13] = soc1.lsu.stq_13_valid;
	assign stq_valids_1[14] = soc1.lsu.stq_14_valid;
	assign stq_valids_1[15] = soc1.lsu.stq_15_valid;

	wire lcam_stq_idx_valid_1;
	assign lcam_stq_idx_valid_1 = 
	//if a load got fired, its stq entry has to be valid
	(soc1.lsu.fired_sta_incoming_REG || soc1.lsu.fired_stad_incoming_REG || soc1.lsu.fired_sta_retry_REG) && !soc1.lsu.REG_1 ? stq_valids_1[soc1.lsu.lcam_stq_idx_0] : 1'b1;
	
	wire ldq_consistent_rob_idx_1;
	assign ldq_consistent_rob_idx_1 =
	  (ldq_valids_1[soc1.lsu.ldq_head])
	  ?
	    (ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 0) % 16], soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx) ? 1'b1 : (soc1.core.rob.full && (soc1.core.rob.io_rob_head_idx == soc1.core.rob.io_rob_tail_idx))) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 1) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 0) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 1) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 2) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 1) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 2) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 3) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 2) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 3) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 4) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 3) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 4) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 5) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 4) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 5) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 6) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 5) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 6) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 7) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 6) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 7) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 8) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 7) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 8) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 9) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 8) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 9) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 10) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 9) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 10) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 11) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 10) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 11) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 12) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 11) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 12) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 13) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 12) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 13) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 14) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 13) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 14) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_1[(soc1.lsu.ldq_head + 15) % 16] ? ROBisOlder(ldq_rob_idx_1[(soc1.lsu.ldq_head + 14) % 16], ldq_rob_idx_1[(soc1.lsu.ldq_head + 15) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1)
	  :
	  	1'b1;

	wire stq_consistent_rob_idx_1;
	assign stq_consistent_rob_idx_1 =
	  stq_valids_1[soc1.lsu.stq_head]
		  ?
	    (ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 0) % 16], soc1.core.rob.io_rob_tail_idx, soc1.core.rob.io_rob_head_idx) ? 1'b1 : (stq_committed_1[(soc1.lsu.stq_head + 0) % 16]) || (soc1.core.rob.full && (soc1.core.rob.io_rob_head_idx == soc1.core.rob.io_rob_tail_idx))) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 1) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 1) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 0) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 0) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 1) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 2) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 2) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 1) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 1) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 2) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 3) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 3) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 2) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 2) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 3) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 4) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 4) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 3) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 3) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 4) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 5) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 5) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 4) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 4) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 5) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 6) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 6) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 5) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 5) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 6) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 7) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 7) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 6) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 6) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 7) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 8) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 8) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 7) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 7) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 8) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 9) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 9) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 8) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 8) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 9) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 10) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 10) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 9) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 9) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 10) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 11) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 11) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 10) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 10) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 11) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 12) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 12) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 11) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 11) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 12) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 13) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 13) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 12) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 12) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 13) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 14) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 14) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 13) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 13) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 14) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_1[(soc1.lsu.stq_head + 15) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 15) % 16] && !stq_committed_1[(soc1.lsu.stq_head + 14) % 16] ? ROBisOlder(stq_rob_idx_1[(soc1.lsu.stq_head + 14) % 16], stq_rob_idx_1[(soc1.lsu.stq_head + 15) % 16], soc1.core.rob.io_rob_head_idx) : 1'b1)
	  :
	  	1'b1;
	
	wire consistent_stq_committed_1;
	assign consistent_stq_committed_1 =
	(soc1.lsu.stq_0_bits_committed ? soc1.lsu.stq_0_valid : 1'b1) &&
	(soc1.lsu.stq_1_bits_committed ? soc1.lsu.stq_1_valid : 1'b1) &&
	(soc1.lsu.stq_2_bits_committed ? soc1.lsu.stq_2_valid : 1'b1) &&
	(soc1.lsu.stq_3_bits_committed ? soc1.lsu.stq_3_valid : 1'b1) &&
	(soc1.lsu.stq_4_bits_committed ? soc1.lsu.stq_4_valid : 1'b1) &&
	(soc1.lsu.stq_5_bits_committed ? soc1.lsu.stq_5_valid : 1'b1) &&
	(soc1.lsu.stq_6_bits_committed ? soc1.lsu.stq_6_valid : 1'b1) &&
	(soc1.lsu.stq_7_bits_committed ? soc1.lsu.stq_7_valid : 1'b1) &&
	(soc1.lsu.stq_8_bits_committed ? soc1.lsu.stq_8_valid : 1'b1) &&
	(soc1.lsu.stq_9_bits_committed ? soc1.lsu.stq_9_valid : 1'b1) &&
	(soc1.lsu.stq_10_bits_committed ? soc1.lsu.stq_10_valid : 1'b1) &&
	(soc1.lsu.stq_11_bits_committed ? soc1.lsu.stq_11_valid : 1'b1) &&
	(soc1.lsu.stq_12_bits_committed ? soc1.lsu.stq_12_valid : 1'b1) &&
	(soc1.lsu.stq_13_bits_committed ? soc1.lsu.stq_13_valid : 1'b1) &&
	(soc1.lsu.stq_14_bits_committed ? soc1.lsu.stq_14_valid : 1'b1) &&
	(soc1.lsu.stq_15_bits_committed ? soc1.lsu.stq_15_valid : 1'b1);	
	
	wire committed_stores_not_speculative_1;
	assign committed_stores_not_speculative_1 =
	  (soc1.lsu.stq_0_bits_committed ? soc1.lsu.stq_0_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_1_bits_committed ? soc1.lsu.stq_1_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_2_bits_committed ? soc1.lsu.stq_2_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_3_bits_committed ? soc1.lsu.stq_3_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_4_bits_committed ? soc1.lsu.stq_4_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_5_bits_committed ? soc1.lsu.stq_5_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_6_bits_committed ? soc1.lsu.stq_6_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_7_bits_committed ? soc1.lsu.stq_7_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_8_bits_committed ? soc1.lsu.stq_8_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_9_bits_committed ? soc1.lsu.stq_9_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_10_bits_committed ? soc1.lsu.stq_10_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_11_bits_committed ? soc1.lsu.stq_11_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_12_bits_committed ? soc1.lsu.stq_12_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_13_bits_committed ? soc1.lsu.stq_13_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_14_bits_committed ? soc1.lsu.stq_14_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.lsu.stq_15_bits_committed ? soc1.lsu.stq_15_bits_uop_br_mask == 12'b0 : 1'b1);
	  
  	wire ldq_rob_valid_consistency_1;
	assign ldq_rob_valid_consistency_1 =
	  (soc1.lsu.ldq_0_valid ? rob_valids_1[soc1.lsu.ldq_0_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_1_valid ? rob_valids_1[soc1.lsu.ldq_1_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_2_valid ? rob_valids_1[soc1.lsu.ldq_2_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_3_valid ? rob_valids_1[soc1.lsu.ldq_3_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_4_valid ? rob_valids_1[soc1.lsu.ldq_4_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_5_valid ? rob_valids_1[soc1.lsu.ldq_5_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_6_valid ? rob_valids_1[soc1.lsu.ldq_6_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_7_valid ? rob_valids_1[soc1.lsu.ldq_7_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_8_valid ? rob_valids_1[soc1.lsu.ldq_8_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_9_valid ? rob_valids_1[soc1.lsu.ldq_9_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_10_valid ? rob_valids_1[soc1.lsu.ldq_10_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_11_valid ? rob_valids_1[soc1.lsu.ldq_11_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_12_valid ? rob_valids_1[soc1.lsu.ldq_12_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_13_valid ? rob_valids_1[soc1.lsu.ldq_13_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_14_valid ? rob_valids_1[soc1.lsu.ldq_14_bits_uop_rob_idx] : 1'b1) &&
	  (soc1.lsu.ldq_15_valid ? rob_valids_1[soc1.lsu.ldq_15_bits_uop_rob_idx] : 1'b1);

	wire speculative_store_rpq_1;
	assign speculative_store_rpq_1 =
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_0 && soc1.dcache.mshrs.mshrs_0.rpq.uops_0_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_1 && soc1.dcache.mshrs.mshrs_0.rpq.uops_1_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_2 && soc1.dcache.mshrs.mshrs_0.rpq.uops_2_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_3 && soc1.dcache.mshrs.mshrs_0.rpq.uops_3_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_4 && soc1.dcache.mshrs.mshrs_0.rpq.uops_4_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_5 && soc1.dcache.mshrs.mshrs_0.rpq.uops_5_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_6 && soc1.dcache.mshrs.mshrs_0.rpq.uops_6_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_7 && soc1.dcache.mshrs.mshrs_0.rpq.uops_7_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_8 && soc1.dcache.mshrs.mshrs_0.rpq.uops_8_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_9 && soc1.dcache.mshrs.mshrs_0.rpq.uops_9_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_10 && soc1.dcache.mshrs.mshrs_0.rpq.uops_10_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_11 && soc1.dcache.mshrs.mshrs_0.rpq.uops_11_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_12 && soc1.dcache.mshrs.mshrs_0.rpq.uops_12_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_13 && soc1.dcache.mshrs.mshrs_0.rpq.uops_13_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_14 && soc1.dcache.mshrs.mshrs_0.rpq.uops_14_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_0.rpq.valids_15 && soc1.dcache.mshrs.mshrs_0.rpq.uops_15_uses_stq && (soc1.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_0 && soc1.dcache.mshrs.mshrs_1.rpq.uops_0_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_1 && soc1.dcache.mshrs.mshrs_1.rpq.uops_1_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_2 && soc1.dcache.mshrs.mshrs_1.rpq.uops_2_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_3 && soc1.dcache.mshrs.mshrs_1.rpq.uops_3_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_4 && soc1.dcache.mshrs.mshrs_1.rpq.uops_4_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_5 && soc1.dcache.mshrs.mshrs_1.rpq.uops_5_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_6 && soc1.dcache.mshrs.mshrs_1.rpq.uops_6_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_7 && soc1.dcache.mshrs.mshrs_1.rpq.uops_7_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_8 && soc1.dcache.mshrs.mshrs_1.rpq.uops_8_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_9 && soc1.dcache.mshrs.mshrs_1.rpq.uops_9_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_10 && soc1.dcache.mshrs.mshrs_1.rpq.uops_10_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_11 && soc1.dcache.mshrs.mshrs_1.rpq.uops_11_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_12 && soc1.dcache.mshrs.mshrs_1.rpq.uops_12_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_13 && soc1.dcache.mshrs.mshrs_1.rpq.uops_13_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_14 && soc1.dcache.mshrs.mshrs_1.rpq.uops_14_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask != 12'b0)) ||
	  (soc1.dcache.mshrs.mshrs_1.rpq.valids_15 && soc1.dcache.mshrs.mshrs_1.rpq.uops_15_uses_stq && (soc1.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask != 12'b0));
	
	wire speculative_store_s1_s2_1;
	assign speculative_store_s1_s2_1 =
	  (soc1.dcache.s1_valid_REG && soc1.dcache.s1_req_0_uop_uses_stq ? soc1.dcache.s1_req_0_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc1.dcache.s2_valid_REG && soc1.dcache.s2_req_0_uop_uses_stq ? soc1.dcache.s2_req_0_uop_br_mask == 12'b0 : 1'b1);
	  
	  
	wire fpiu_BranchKillableQueue_1_not_committed_1;
	assign fpiu_BranchKillableQueue_1_not_committed_1 =
	  (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0 ? !(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_stq_idx]) : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1 ? !(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_stq_idx]) : 1'b1) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2 ? !(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_uses_stq && stq_committed_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_stq_idx]) : 1'b1);

	wire fdivsqrt_valid_consistency_1;
	assign fdivsqrt_valid_consistency_1 = soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.io_outValid_div || soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.io_outValid_sqrt ? soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val : 1'b1;

	wire div_state_1;
	assign div_state_1 = !soc1.core.reset ? (soc1.core.csr_exe_unit.div.div.state == 3'h0) || (soc1.core.csr_exe_unit.div.div.state == 3'h3) || (soc1.core.csr_exe_unit.div.div.state == 3'h7) : 1'b1;

	wire ldq_entries_not_using_stq_1;
	assign ldq_entries_not_using_stq_1 = 
	  !soc1.lsu.ldq_0_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_1_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_2_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_3_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_4_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_5_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_6_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_7_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_8_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_9_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_10_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_11_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_12_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_13_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_14_bits_uop_uses_stq &&
	  !soc1.lsu.ldq_15_bits_uop_uses_stq;

	wire stq_entries_not_using_ldq_1;
	assign stq_entries_not_using_ldq_1 = 
	  !soc1.lsu.stq_0_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_1_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_2_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_3_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_4_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_5_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_6_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_7_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_8_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_9_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_10_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_11_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_12_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_13_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_14_bits_uop_uses_ldq &&
	  !soc1.lsu.stq_15_bits_uop_uses_ldq;
	  
	wire BranchKillableQueue_empty_1;
	assign BranchKillableQueue_empty_1 =
	soc1.core.b2_mispredict ||
	(soc1.core.jmp_unit.queue.io_empty ==
	(!soc1.core.jmp_unit.queue.valids_0 &&
	!soc1.core.jmp_unit.queue.valids_1 &&
	!soc1.core.jmp_unit.queue.valids_2 &&
	!soc1.core.jmp_unit.queue.valids_3 &&
	!soc1.core.jmp_unit.queue.valids_4)) &&

	(soc1.core.fp_pipeline.fpiu_unit.queue.io_empty ==
	(!soc1.core.fp_pipeline.fpiu_unit.queue.valids_0 &&
	!soc1.core.fp_pipeline.fpiu_unit.queue.valids_1 &&
	!soc1.core.fp_pipeline.fpiu_unit.queue.valids_2 &&
	!soc1.core.fp_pipeline.fpiu_unit.queue.valids_3 &&
	!soc1.core.fp_pipeline.fpiu_unit.queue.valids_4 &&
	!soc1.core.fp_pipeline.fpiu_unit.queue.valids_5 &&
	!soc1.core.fp_pipeline.fpiu_unit.queue.valids_6)) &&

	(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.io_empty ==
	(!soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0 &&
	!soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1 &&
	!soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2)) &&

	(
	  (soc1.core.jmp_unit.queue.value == 3'h0 && soc1.core.jmp_unit.queue.valids_0) ||
	  (soc1.core.jmp_unit.queue.value == 3'h1 && soc1.core.jmp_unit.queue.valids_1) ||
	  (soc1.core.jmp_unit.queue.value == 3'h2 && soc1.core.jmp_unit.queue.valids_2) ||
	  (soc1.core.jmp_unit.queue.value == 3'h3 && soc1.core.jmp_unit.queue.valids_3) ||
	  (soc1.core.jmp_unit.queue.value == 3'h4 && soc1.core.jmp_unit.queue.valids_4)
	  ?
	  !soc1.core.jmp_unit.queue.do_enq
	  :
	  1'b1
	) &&
	(
	  (soc1.core.fp_pipeline.fpiu_unit.queue.value == 3'h0 && soc1.core.fp_pipeline.fpiu_unit.queue.valids_0) ||
	  (soc1.core.fp_pipeline.fpiu_unit.queue.value == 3'h1 && soc1.core.fp_pipeline.fpiu_unit.queue.valids_1) ||
	  (soc1.core.fp_pipeline.fpiu_unit.queue.value == 3'h2 && soc1.core.fp_pipeline.fpiu_unit.queue.valids_2) ||
	  (soc1.core.fp_pipeline.fpiu_unit.queue.value == 3'h3 && soc1.core.fp_pipeline.fpiu_unit.queue.valids_3) ||
	  (soc1.core.fp_pipeline.fpiu_unit.queue.value == 3'h4 && soc1.core.fp_pipeline.fpiu_unit.queue.valids_4) ||
	  (soc1.core.fp_pipeline.fpiu_unit.queue.value == 3'h5 && soc1.core.fp_pipeline.fpiu_unit.queue.valids_5) ||
	  (soc1.core.fp_pipeline.fpiu_unit.queue.value == 3'h6 && soc1.core.fp_pipeline.fpiu_unit.queue.valids_6)
	  ?
	  !soc1.core.fp_pipeline.fpiu_unit.queue.do_enq
	  :
	  1'b1
	) &&
	(
	  (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value == 2'h0 && soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0) ||
	  (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value == 2'h1 && soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1) ||
	  (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value == 2'h2 && soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2)
	  ?
	  !soc1.core.fp_pipeline.fpiu_unit.fp_sdq.do_enq
	  :
	  1'b1
	);
	
		
	wire BranchKillableQueue_pointers_valid_1;
	assign BranchKillableQueue_pointers_valid_1 =
	(soc1.core.jmp_unit.queue.value < 3'h5) && (soc1.core.jmp_unit.queue.value_1 < 3'h5) &&
	(soc1.core.fp_pipeline.fpiu_unit.queue.value < 3'h7) && (soc1.core.fp_pipeline.fpiu_unit.queue.value_1 < 3'h7) &&
	(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value < 2'h3) && (soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 < 2'h3)
	;
	
	wire [5:0] bkq_jmp_rob_idx_1 [4:0];
	assign bkq_jmp_rob_idx_1[0] = soc1.core.jmp_unit.queue.uops_0_rob_idx;
	assign bkq_jmp_rob_idx_1[1] = soc1.core.jmp_unit.queue.uops_1_rob_idx;
	assign bkq_jmp_rob_idx_1[2] = soc1.core.jmp_unit.queue.uops_2_rob_idx;
	assign bkq_jmp_rob_idx_1[3] = soc1.core.jmp_unit.queue.uops_3_rob_idx;
	assign bkq_jmp_rob_idx_1[4] = soc1.core.jmp_unit.queue.uops_4_rob_idx;

	wire bkq_jmp_valids_1 [4:0];
	assign bkq_jmp_valids_1[0] = soc1.core.jmp_unit.queue.valids_0;
	assign bkq_jmp_valids_1[1] = soc1.core.jmp_unit.queue.valids_1;
	assign bkq_jmp_valids_1[2] = soc1.core.jmp_unit.queue.valids_2;
	assign bkq_jmp_valids_1[3] = soc1.core.jmp_unit.queue.valids_3;
	assign bkq_jmp_valids_1[4] = soc1.core.jmp_unit.queue.valids_4;
	  
	wire bkq_jmp_rob_consistency_1;
	assign bkq_jmp_rob_consistency_1 =
	!soc1.core.jmp_unit.queue.io_empty
	?
	  (bkq_jmp_valids_1[(soc1.core.jmp_unit.queue.value_1 + 1) % 5] ? ROBisOlder(bkq_jmp_rob_idx_1[soc1.core.jmp_unit.queue.value_1], bkq_jmp_rob_idx_1[(soc1.core.jmp_unit.queue.value_1 + 1) % 5], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_jmp_valids_1[(soc1.core.jmp_unit.queue.value_1 + 2) % 5] ? ROBisOlder(bkq_jmp_rob_idx_1[(soc1.core.jmp_unit.queue.value_1 + 1) % 5], bkq_jmp_rob_idx_1[(soc1.core.jmp_unit.queue.value_1 + 2) % 5], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_jmp_valids_1[(soc1.core.jmp_unit.queue.value_1 + 3) % 5] ? ROBisOlder(bkq_jmp_rob_idx_1[(soc1.core.jmp_unit.queue.value_1 + 2) % 5], bkq_jmp_rob_idx_1[(soc1.core.jmp_unit.queue.value_1 + 3) % 5], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_jmp_valids_1[(soc1.core.jmp_unit.queue.value_1 + 4) % 5] ? ROBisOlder(bkq_jmp_rob_idx_1[(soc1.core.jmp_unit.queue.value_1 + 3) % 5], bkq_jmp_rob_idx_1[(soc1.core.jmp_unit.queue.value_1 + 4) % 5], soc1.core.rob.io_rob_head_idx) : 1'b1)
	:
	  1'b1;

	wire [5:0] bkq_fp_rob_idx_1 [6:0];
	assign bkq_fp_rob_idx_1[0] = soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx;
	assign bkq_fp_rob_idx_1[1] = soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx;
	assign bkq_fp_rob_idx_1[2] = soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx;
	assign bkq_fp_rob_idx_1[3] = soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx;
	assign bkq_fp_rob_idx_1[4] = soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx;
	assign bkq_fp_rob_idx_1[5] = soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx;
	assign bkq_fp_rob_idx_1[6] = soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx;


	wire bkq_fp_valids_1 [6:0];
	assign bkq_fp_valids_1[0] = soc1.core.fp_pipeline.fpiu_unit.queue.valids_0;
	assign bkq_fp_valids_1[1] = soc1.core.fp_pipeline.fpiu_unit.queue.valids_1;
	assign bkq_fp_valids_1[2] = soc1.core.fp_pipeline.fpiu_unit.queue.valids_2;
	assign bkq_fp_valids_1[3] = soc1.core.fp_pipeline.fpiu_unit.queue.valids_3;
	assign bkq_fp_valids_1[4] = soc1.core.fp_pipeline.fpiu_unit.queue.valids_4;
	assign bkq_fp_valids_1[5] = soc1.core.fp_pipeline.fpiu_unit.queue.valids_5;
	assign bkq_fp_valids_1[6] = soc1.core.fp_pipeline.fpiu_unit.queue.valids_6;

	wire bkq_fp_rob_consistency_1;
	assign bkq_fp_rob_consistency_1 =
	!soc1.core.fp_pipeline.fpiu_unit.queue.io_empty
	?
	  (bkq_fp_valids_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 1) % 7] ? ROBisOlder(bkq_fp_rob_idx_1[soc1.core.fp_pipeline.fpiu_unit.queue.value_1], bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 1) % 7], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 2) % 7] ? ROBisOlder(bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 1) % 7], bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 2) % 7], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 3) % 7] ? ROBisOlder(bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 2) % 7], bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 3) % 7], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 4) % 7] ? ROBisOlder(bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 3) % 7], bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 4) % 7], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 5) % 7] ? ROBisOlder(bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 4) % 7], bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 5) % 7], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 6) % 7] ? ROBisOlder(bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 5) % 7], bkq_fp_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.queue.value_1 + 6) % 7], soc1.core.rob.io_rob_head_idx) : 1'b1)
	:
	  1'b1;

	wire [5:0] bkq_fp_1_rob_idx_1 [2:0];
	assign bkq_fp_1_rob_idx_1[0] = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx;
	assign bkq_fp_1_rob_idx_1[1] = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx;
	assign bkq_fp_1_rob_idx_1[2] = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx;

	wire bkq_fp_1_valids_1 [2:0];
	assign bkq_fp_1_valids_1[0] = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0;
	assign bkq_fp_1_valids_1[1] = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1;
	assign bkq_fp_1_valids_1[2] = soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2;
	  
	wire bkq_fp_1_rob_consistency_1;
	assign bkq_fp_1_rob_consistency_1 =
	!soc1.core.fp_pipeline.fpiu_unit.fp_sdq.io_empty
	?
	  (bkq_fp_1_valids_1[(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 1) % 3] ? ROBisOlder(bkq_fp_1_rob_idx_1[soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value_1], bkq_fp_1_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 1) % 3], soc1.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_1_valids_1[(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 2) % 3] ? ROBisOlder(bkq_fp_1_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 1) % 3], bkq_fp_1_rob_idx_1[(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 2) % 3], soc1.core.rob.io_rob_head_idx) : 1'b1)
	:
	  1'b1;

	/*wire ROB_uops_equal_STQ_1;
	assign ROB_uops_equal_STQ_1 =
	  ROB_exists_in_STQ(6'h0, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h1, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h2, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h3, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h4, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h5, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h6, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h7, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h8, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h9, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'ha, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'hb, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'hc, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'hd, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'he, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'hf, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h10, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h11, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h12, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h13, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h14, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h15, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h16, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h17, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h18, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h19, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h1a, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h1b, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h1c, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h1d, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h1e, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h1f, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h20, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h21, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h22, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h23, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h24, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h25, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h26, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h27, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h28, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h29, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h2a, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h2b, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h2c, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h2d, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h2e, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h2f, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h30, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h31, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h32, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h33, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h34, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h35, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h36, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h37, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h38, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h39, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h3a, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h3b, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h3c, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h3d, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h3e, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1) &&
	  ROB_exists_in_STQ(6'h3f, rob_valids_1, rob_uses_stq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, stq_rob_idx_1, rob_stq_indexes_1, stq_valids_1, stq_committed_1);

	wire ROB_uops_equal_LDQ_1;
	assign ROB_uops_equal_LDQ_1 =
	  ROB_exists_in_LDQ(6'h0, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h1, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h2, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h3, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h4, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h5, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h6, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h7, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h8, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h9, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'ha, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'hb, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'hc, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'hd, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'he, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'hf, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h10, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h11, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h12, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h13, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h14, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h15, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h16, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h17, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h18, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h19, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h1a, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h1b, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h1c, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h1d, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h1e, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h1f, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h20, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h21, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h22, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h23, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h24, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h25, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h26, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h27, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h28, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h29, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h2a, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h2b, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h2c, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h2d, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h2e, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h2f, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h30, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h31, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h32, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h33, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h34, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h35, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h36, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h37, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h38, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h39, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h3a, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h3b, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h3c, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h3d, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h3e, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1) &&
	  ROB_exists_in_LDQ(6'h3f, rob_valids_1, rob_uses_ldq_1, soc1.core.rob.rob_state, soc1.core.rob.REG_1, rob_exception_1, ldq_rob_idx_1, rob_ldq_indexes_1, ldq_valids_1);*/

	wire STQ_uops_equals_ROB_1;
	assign STQ_uops_equals_ROB_1 =
	  STQ_exists_in_ROB(4'h0, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'h1, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'h2, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'h3, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'h4, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'h5, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'h6, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'h7, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'h8, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'h9, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'ha, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'hb, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'hc, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'hd, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'he, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1) &&
	  STQ_exists_in_ROB(4'hf, stq_valids_1, stq_committed_1, rob_uses_stq_1, stq_rob_idx_1, rob_valids_1);

	wire LDQ_uops_equals_ROB_1;
	assign LDQ_uops_equals_ROB_1 =
	  LDQ_exists_in_ROB(4'h0, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'h1, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'h2, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'h3, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'h4, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'h5, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'h6, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'h7, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'h8, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'h9, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'ha, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'hb, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'hc, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'hd, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'he, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1) &&
	  LDQ_exists_in_ROB(4'hf, ldq_valids_1, rob_uses_ldq_1, ldq_rob_idx_1, rob_valids_1);
	  
	wire ldq_uses_ldq_1[15:0];
	assign ldq_uses_ldq_1[0] = soc1.lsu.ldq_0_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[1] = soc1.lsu.ldq_1_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[2] = soc1.lsu.ldq_2_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[3] = soc1.lsu.ldq_3_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[4] = soc1.lsu.ldq_4_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[5] = soc1.lsu.ldq_5_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[6] = soc1.lsu.ldq_6_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[7] = soc1.lsu.ldq_7_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[8] = soc1.lsu.ldq_8_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[9] = soc1.lsu.ldq_9_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[10] = soc1.lsu.ldq_10_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[11] = soc1.lsu.ldq_11_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[12] = soc1.lsu.ldq_12_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[13] = soc1.lsu.ldq_13_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[14] = soc1.lsu.ldq_14_bits_uop_uses_ldq;
	assign ldq_uses_ldq_1[15] = soc1.lsu.ldq_15_bits_uop_uses_ldq;
	  
	wire stq_uses_stq_1[15:0];
	assign stq_uses_stq_1[0] = soc1.lsu.stq_0_bits_uop_uses_stq;
	assign stq_uses_stq_1[1] = soc1.lsu.stq_1_bits_uop_uses_stq;
	assign stq_uses_stq_1[2] = soc1.lsu.stq_2_bits_uop_uses_stq;
	assign stq_uses_stq_1[3] = soc1.lsu.stq_3_bits_uop_uses_stq;
	assign stq_uses_stq_1[4] = soc1.lsu.stq_4_bits_uop_uses_stq;
	assign stq_uses_stq_1[5] = soc1.lsu.stq_5_bits_uop_uses_stq;
	assign stq_uses_stq_1[6] = soc1.lsu.stq_6_bits_uop_uses_stq;
	assign stq_uses_stq_1[7] = soc1.lsu.stq_7_bits_uop_uses_stq;
	assign stq_uses_stq_1[8] = soc1.lsu.stq_8_bits_uop_uses_stq;
	assign stq_uses_stq_1[9] = soc1.lsu.stq_9_bits_uop_uses_stq;
	assign stq_uses_stq_1[10] = soc1.lsu.stq_10_bits_uop_uses_stq;
	assign stq_uses_stq_1[11] = soc1.lsu.stq_11_bits_uop_uses_stq;
	assign stq_uses_stq_1[12] = soc1.lsu.stq_12_bits_uop_uses_stq;
	assign stq_uses_stq_1[13] = soc1.lsu.stq_13_bits_uop_uses_stq;
	assign stq_uses_stq_1[14] = soc1.lsu.stq_14_bits_uop_uses_stq;
	assign stq_uses_stq_1[15] = soc1.lsu.stq_15_bits_uop_uses_stq;
	  
	wire buffers_equal_ROB_1;
	assign buffers_equal_ROB_1 =
	Buffer_exists_in_ROB_stq_idx_only(soc1.core.b2_mispredict, stq_committed_1, soc1.core.b2_uop_stq_idx, rob_valids_1, soc1.core.b2_uop_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc1.core.brinfos_0_valid, stq_committed_1, soc1.core.brinfos_0_uop_stq_idx, rob_valids_1, soc1.core.brinfos_0_uop_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc1.core.brinfos_1_valid, stq_committed_1, soc1.core.brinfos_1_uop_stq_idx, rob_valids_1, soc1.core.brinfos_1_uop_rob_idx) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.csr_exe_unit.alu.r_valids_0, soc1.core.csr_exe_unit.alu.r_uops_0_uses_stq, rob_valids_1, soc1.core.csr_exe_unit.alu.r_uops_0_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq((soc1.core.csr_exe_unit.div.div.state == 3'h3) || (soc1.core.csr_exe_unit.div.div.state == 3'h7), soc1.core.csr_exe_unit.div.r_uop_uses_stq, rob_valids_1, soc1.core.csr_exe_unit.div.r_uop_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_0.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_1.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_2.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_3.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_4.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_5.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_6.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_7.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_8.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_9.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_10.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_11.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_12.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_13.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_14.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fp_issue_unit.slots_15.io_valid, soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.queue.valids_0, soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.queue.valids_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.queue.valids_2, soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.queue.valids_3, soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.queue.valids_4, soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.queue.valids_5, soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.queue.valids_6, soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_no_idx(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_val, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_uses_stq, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_uses_ldq) &&
	Buffer_exists_in_ROB_no_idx(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_uses_stq, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_uses_ldq) &&
	Buffer_exists_in_ROB_no_idx(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_val, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_uses_stq, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_0, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_2, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fpiu_unit.fpu.r_valids_3, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fregister_read.exe_reg_valids_0, soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx, rob_uses_stq_1, rob_uses_ldq_1,soc1.core.fp_pipeline.fregister_read.exe_reg_uops_0_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.fp_pipeline.fregister_read.rrd_valids_0_REG, soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uses_stq, stq_committed_1, soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_stq_idx, rob_valids_1, soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx, rob_uses_stq_1, rob_uses_ldq_1,soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_0.io_valid, soc1.core.int_issue_unit.slots_0.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_0.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_0.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_0.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_1.io_valid, soc1.core.int_issue_unit.slots_1.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_1.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_1.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_1.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_2.io_valid, soc1.core.int_issue_unit.slots_2.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_2.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_2.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_2.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_3.io_valid, soc1.core.int_issue_unit.slots_3.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_3.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_3.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_3.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_4.io_valid, soc1.core.int_issue_unit.slots_4.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_4.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_4.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_4.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_5.io_valid, soc1.core.int_issue_unit.slots_5.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_5.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_5.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_5.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_6.io_valid, soc1.core.int_issue_unit.slots_6.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_6.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_6.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_6.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_7.io_valid, soc1.core.int_issue_unit.slots_7.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_7.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_7.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_7.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_8.io_valid, soc1.core.int_issue_unit.slots_8.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_8.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_8.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_8.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_9.io_valid, soc1.core.int_issue_unit.slots_9.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_9.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_9.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_9.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_10.io_valid, soc1.core.int_issue_unit.slots_10.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_10.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_10.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_10.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_11.io_valid, soc1.core.int_issue_unit.slots_11.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_11.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_11.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_11.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_12.io_valid, soc1.core.int_issue_unit.slots_12.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_12.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_12.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_12.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_13.io_valid, soc1.core.int_issue_unit.slots_13.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_13.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_13.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_13.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_14.io_valid, soc1.core.int_issue_unit.slots_14.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_14.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_14.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_14.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_15.io_valid, soc1.core.int_issue_unit.slots_15.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_15.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_15.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_15.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_16.io_valid, soc1.core.int_issue_unit.slots_16.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_16.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_16.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_16.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_17.io_valid, soc1.core.int_issue_unit.slots_17.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_17.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_17.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_17.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_18.io_valid, soc1.core.int_issue_unit.slots_18.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_18.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_18.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_18.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.int_issue_unit.slots_19.io_valid, soc1.core.int_issue_unit.slots_19.slot_uop_uses_stq, stq_committed_1, soc1.core.int_issue_unit.slots_19.slot_uop_stq_idx, rob_valids_1, soc1.core.int_issue_unit.slots_19.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.int_issue_unit.slots_19.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.iregister_read.exe_reg_valids_0, soc1.core.iregister_read.exe_reg_uops_0_uses_stq, stq_committed_1, soc1.core.iregister_read.exe_reg_uops_0_stq_idx, rob_valids_1, soc1.core.iregister_read.exe_reg_uops_0_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.iregister_read.exe_reg_uops_0_uses_ldq) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.iregister_read.exe_reg_valids_1, soc1.core.iregister_read.exe_reg_uops_1_uses_stq, stq_committed_1, soc1.core.iregister_read.exe_reg_uops_1_stq_idx, rob_valids_1, soc1.core.iregister_read.exe_reg_uops_1_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.iregister_read.exe_reg_valids_2, soc1.core.iregister_read.exe_reg_uops_2_uses_stq, stq_committed_1, soc1.core.iregister_read.exe_reg_uops_2_stq_idx, rob_valids_1, soc1.core.iregister_read.exe_reg_uops_2_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB(soc1.core.iregister_read.rrd_valids_0_REG, soc1.core.iregister_read.rrd_uops_0_REG_uses_stq, stq_committed_1, soc1.core.iregister_read.rrd_uops_0_REG_stq_idx, rob_valids_1, soc1.core.iregister_read.rrd_uops_0_REG_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.iregister_read.rrd_uops_0_REG_uses_ldq) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.iregister_read.rrd_valids_1_REG, soc1.core.iregister_read.rrd_uops_1_REG_uses_stq, stq_committed_1, soc1.core.iregister_read.rrd_uops_1_REG_stq_idx, rob_valids_1, soc1.core.iregister_read.rrd_uops_1_REG_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_stq(soc1.core.iregister_read.rrd_valids_2_REG, soc1.core.iregister_read.rrd_uops_2_REG_uses_stq, stq_committed_1, soc1.core.iregister_read.rrd_uops_2_REG_stq_idx, rob_valids_1, soc1.core.iregister_read.rrd_uops_2_REG_rob_idx, rob_uses_stq_1) &&
	//(soc1.core.jmp_unit.queue.ram_fflags_valid ? rob_valids_1[soc1.core.jmp_unit.queue.ram_fflags_bits_uop_rob_idx] : 1'b1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.queue.valids_0, soc1.core.jmp_unit.queue.uops_0_uses_stq, rob_valids_1, soc1.core.jmp_unit.queue.uops_0_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.queue.valids_1, soc1.core.jmp_unit.queue.uops_1_uses_stq, rob_valids_1, soc1.core.jmp_unit.queue.uops_1_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.queue.valids_2, soc1.core.jmp_unit.queue.uops_2_uses_stq, rob_valids_1, soc1.core.jmp_unit.queue.uops_2_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.queue.valids_3, soc1.core.jmp_unit.queue.uops_3_uses_stq, rob_valids_1, soc1.core.jmp_unit.queue.uops_3_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.queue.valids_4, soc1.core.jmp_unit.queue.uops_4_uses_stq, rob_valids_1, soc1.core.jmp_unit.queue.uops_4_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.alu.r_valids_0, soc1.core.jmp_unit.alu.r_uops_0_uses_stq, rob_valids_1, soc1.core.jmp_unit.alu.r_uops_0_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.alu.r_valids_1, soc1.core.jmp_unit.alu.r_uops_1_uses_stq, rob_valids_1, soc1.core.jmp_unit.alu.r_uops_1_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.alu.r_valids_2, soc1.core.jmp_unit.alu.r_uops_2_uses_stq, rob_valids_1, soc1.core.jmp_unit.alu.r_uops_2_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.ifpu.r_valids_0, soc1.core.jmp_unit.ifpu.r_uops_0_uses_stq, rob_valids_1, soc1.core.jmp_unit.ifpu.r_uops_0_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.ifpu.r_valids_1, soc1.core.jmp_unit.ifpu.r_uops_1_uses_stq, rob_valids_1, soc1.core.jmp_unit.ifpu.r_uops_1_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.imul.r_valids_0, soc1.core.jmp_unit.imul.r_uops_0_uses_stq, rob_valids_1, soc1.core.jmp_unit.imul.r_uops_0_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.imul.r_valids_1, soc1.core.jmp_unit.imul.r_uops_1_uses_stq, rob_valids_1, soc1.core.jmp_unit.imul.r_uops_1_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc1.core.jmp_unit.imul.r_valids_2, soc1.core.jmp_unit.imul.r_uops_2_uses_stq, rob_valids_1, soc1.core.jmp_unit.imul.r_uops_2_rob_idx, rob_uses_stq_1) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_0.io_valid, soc1.core.mem_issue_unit.slots_0.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_0.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_0.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_0.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_1.io_valid, soc1.core.mem_issue_unit.slots_1.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_1.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_1.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_1.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_2.io_valid, soc1.core.mem_issue_unit.slots_2.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_2.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_2.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_2.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_3.io_valid, soc1.core.mem_issue_unit.slots_3.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_3.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_3.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_3.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_4.io_valid, soc1.core.mem_issue_unit.slots_4.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_4.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_4.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_4.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_5.io_valid, soc1.core.mem_issue_unit.slots_5.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_5.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_5.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_5.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_6.io_valid, soc1.core.mem_issue_unit.slots_6.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_6.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_6.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_6.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_7.io_valid, soc1.core.mem_issue_unit.slots_7.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_7.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_7.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_7.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_8.io_valid, soc1.core.mem_issue_unit.slots_8.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_8.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_8.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_8.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_9.io_valid, soc1.core.mem_issue_unit.slots_9.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_9.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_9.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_9.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_10.io_valid, soc1.core.mem_issue_unit.slots_10.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_10.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_10.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_10.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc1.core.mem_issue_unit.slots_11.io_valid, soc1.core.mem_issue_unit.slots_11.slot_uop_uses_stq, stq_committed_1, soc1.core.mem_issue_unit.slots_11.slot_uop_stq_idx, rob_valids_1, soc1.core.mem_issue_unit.slots_11.slot_uop_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.core.mem_issue_unit.slots_11.slot_uop_uses_ldq) &&
	(soc1.core.rob.r_xcpt_val ? rob_valids_1[soc1.core.rob.r_xcpt_uop_rob_idx] : 1'b1) &&
	//Buffer_exists_in_LDQ(soc1.dcache.s1_valid_0, soc1.dcache.s1_req_0_uop_uses_ldq, ldq_valids_1, soc1.dcache.s1_req_0_uop_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.s1_valid_0 && (soc1.dcache.s1_type != 3'b0 || soc1.dcache.s1_req_0_uop_is_amo), soc1.dcache.s1_req_0_uop_uses_stq, stq_valids_1, soc1.dcache.s1_req_0_uop_stq_idx, stq_uses_stq_1) &&
	//Buffer_exists_in_LDQ(soc1.dcache.s2_valid_0, soc1.dcache.s2_req_0_uop_uses_ldq, ldq_valids_1, soc1.dcache.s2_req_0_uop_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.s2_valid_0 && (soc1.dcache.s2_type != 3'b0 || soc1.dcache.s2_req_0_uop_is_amo), soc1.dcache.s2_req_0_uop_uses_stq, stq_valids_1, soc1.dcache.s2_req_0_uop_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mmios_0.state != 2'b0, soc1.dcache.mshrs.mmios_0.req_uop_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mmios_0.req_uop_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(!soc1.dcache.mshrs.mmios_0.io_req_valid, soc1.dcache.mshrs.mmios_0.req_uop_uses_stq, stq_valids_1, soc1.dcache.mshrs.mmios_0.req_uop_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_0, soc1.dcache.mshrs.mshrs_0.rpq.uops_0_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_0_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_0, soc1.dcache.mshrs.mshrs_0.rpq.uops_0_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_1_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_1_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_1_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_2, soc1.dcache.mshrs.mshrs_0.rpq.uops_2_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_2_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_2, soc1.dcache.mshrs.mshrs_0.rpq.uops_2_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_3, soc1.dcache.mshrs.mshrs_0.rpq.uops_3_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_3_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_3, soc1.dcache.mshrs.mshrs_0.rpq.uops_3_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_4, soc1.dcache.mshrs.mshrs_0.rpq.uops_4_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_4_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_4, soc1.dcache.mshrs.mshrs_0.rpq.uops_4_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_5, soc1.dcache.mshrs.mshrs_0.rpq.uops_5_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_5_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_5, soc1.dcache.mshrs.mshrs_0.rpq.uops_5_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_6, soc1.dcache.mshrs.mshrs_0.rpq.uops_6_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_6_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_6, soc1.dcache.mshrs.mshrs_0.rpq.uops_6_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_7, soc1.dcache.mshrs.mshrs_0.rpq.uops_7_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_7_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_7, soc1.dcache.mshrs.mshrs_0.rpq.uops_7_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_8, soc1.dcache.mshrs.mshrs_0.rpq.uops_8_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_8_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_8, soc1.dcache.mshrs.mshrs_0.rpq.uops_8_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_9, soc1.dcache.mshrs.mshrs_0.rpq.uops_9_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_9_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_9, soc1.dcache.mshrs.mshrs_0.rpq.uops_9_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_10, soc1.dcache.mshrs.mshrs_0.rpq.uops_10_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_10_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_10, soc1.dcache.mshrs.mshrs_0.rpq.uops_10_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_11, soc1.dcache.mshrs.mshrs_0.rpq.uops_11_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_11_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_11, soc1.dcache.mshrs.mshrs_0.rpq.uops_11_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_12, soc1.dcache.mshrs.mshrs_0.rpq.uops_12_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_12_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_12, soc1.dcache.mshrs.mshrs_0.rpq.uops_12_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_13, soc1.dcache.mshrs.mshrs_0.rpq.uops_13_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_13_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_13, soc1.dcache.mshrs.mshrs_0.rpq.uops_13_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_14, soc1.dcache.mshrs.mshrs_0.rpq.uops_14_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_14_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_14, soc1.dcache.mshrs.mshrs_0.rpq.uops_14_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_15, soc1.dcache.mshrs.mshrs_0.rpq.uops_15_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_15_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_0.rpq.valids_15, soc1.dcache.mshrs.mshrs_0.rpq.uops_15_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_0, soc1.dcache.mshrs.mshrs_1.rpq.uops_0_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_0_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_0, soc1.dcache.mshrs.mshrs_1.rpq.uops_0_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_1_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_1_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_1_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_2, soc1.dcache.mshrs.mshrs_1.rpq.uops_2_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_2_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_2, soc1.dcache.mshrs.mshrs_1.rpq.uops_2_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_3, soc1.dcache.mshrs.mshrs_1.rpq.uops_3_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_3_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_3, soc1.dcache.mshrs.mshrs_1.rpq.uops_3_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_4, soc1.dcache.mshrs.mshrs_1.rpq.uops_4_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_4_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_4, soc1.dcache.mshrs.mshrs_1.rpq.uops_4_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_5, soc1.dcache.mshrs.mshrs_1.rpq.uops_5_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_5_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_5, soc1.dcache.mshrs.mshrs_1.rpq.uops_5_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_6, soc1.dcache.mshrs.mshrs_1.rpq.uops_6_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_6_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_6, soc1.dcache.mshrs.mshrs_1.rpq.uops_6_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_7, soc1.dcache.mshrs.mshrs_1.rpq.uops_7_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_7_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_7, soc1.dcache.mshrs.mshrs_1.rpq.uops_7_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_8, soc1.dcache.mshrs.mshrs_1.rpq.uops_8_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_8_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_8, soc1.dcache.mshrs.mshrs_1.rpq.uops_8_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_9, soc1.dcache.mshrs.mshrs_1.rpq.uops_9_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_9_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_9, soc1.dcache.mshrs.mshrs_1.rpq.uops_9_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_10, soc1.dcache.mshrs.mshrs_1.rpq.uops_10_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_10_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_10, soc1.dcache.mshrs.mshrs_1.rpq.uops_10_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_11, soc1.dcache.mshrs.mshrs_1.rpq.uops_11_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_11_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_11, soc1.dcache.mshrs.mshrs_1.rpq.uops_11_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_12, soc1.dcache.mshrs.mshrs_1.rpq.uops_12_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_12_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_12, soc1.dcache.mshrs.mshrs_1.rpq.uops_12_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_13, soc1.dcache.mshrs.mshrs_1.rpq.uops_13_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_13_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_13, soc1.dcache.mshrs.mshrs_1.rpq.uops_13_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_14, soc1.dcache.mshrs.mshrs_1.rpq.uops_14_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_14_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_14, soc1.dcache.mshrs.mshrs_1.rpq.uops_14_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_15, soc1.dcache.mshrs.mshrs_1.rpq.uops_15_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_15_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.mshrs_1.rpq.valids_15, soc1.dcache.mshrs.mshrs_1.rpq.uops_15_uses_stq, stq_valids_1, soc1.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.respq.valids_0, soc1.dcache.mshrs.respq.uops_0_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.respq.uops_0_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.respq.valids_0, soc1.dcache.mshrs.respq.uops_0_uses_stq, stq_valids_1, soc1.dcache.mshrs.respq.uops_0_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.respq.valids_1, soc1.dcache.mshrs.respq.uops_1_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.respq.uops_1_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.respq.valids_1, soc1.dcache.mshrs.respq.uops_1_uses_stq, stq_valids_1, soc1.dcache.mshrs.respq.uops_1_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.respq.valids_2, soc1.dcache.mshrs.respq.uops_2_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.respq.uops_2_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.respq.valids_2, soc1.dcache.mshrs.respq.uops_2_uses_stq, stq_valids_1, soc1.dcache.mshrs.respq.uops_2_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_LDQ(soc1.dcache.mshrs.respq.valids_3, soc1.dcache.mshrs.respq.uops_3_uses_ldq, ldq_valids_1, soc1.dcache.mshrs.respq.uops_3_ldq_idx, ldq_uses_ldq_1) &&
	//Buffer_exists_in_STQ(soc1.dcache.mshrs.respq.valids_3, soc1.dcache.mshrs.respq.uops_3_uses_stq, stq_valids_1, soc1.dcache.mshrs.respq.uops_3_stq_idx, stq_uses_stq_1) &&
	Buffer_exists_in_ROB_stq_idx_only(soc1.lsu.fired_sfence_0 || soc1.lsu.fired_load_incoming_REG || soc1.lsu.fired_sta_incoming_REG || soc1.lsu.fired_stad_incoming_REG || soc1.lsu.fired_std_incoming_REG, stq_committed_1, soc1.lsu.mem_incoming_uop_0_stq_idx, rob_valids_1, soc1.lsu.mem_incoming_uop_0_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc1.lsu.fired_stdf_incoming, stq_committed_1, soc1.lsu.mem_stdf_uop_stq_idx, rob_valids_1, soc1.lsu.mem_stdf_uop_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc1.lsu.fired_sta_incoming_REG || soc1.lsu.fired_stad_incoming_REG || soc1.lsu.fired_std_incoming_REG, stq_committed_1, soc1.lsu.mem_stq_incoming_e_0_bits_uop_stq_idx, rob_valids_1, soc1.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc1.lsu.fired_sta_retry_REG, stq_committed_1, soc1.lsu.mem_stq_retry_e_bits_uop_stq_idx, rob_valids_1, soc1.lsu.mem_stq_retry_e_bits_uop_rob_idx) &&
	Buffer_exists_in_ROB(soc1.lsu.mem_xcpt_valids_0, soc1.lsu.mem_xcpt_uops_0_uses_stq, stq_committed_1, soc1.lsu.mem_xcpt_uops_0_stq_idx, rob_valids_1, soc1.lsu.mem_xcpt_uops_0_rob_idx, rob_uses_stq_1, rob_uses_ldq_1, soc1.lsu.mem_xcpt_uops_0_uses_ldq)
	;
	
	/*function automatic check_uniqueness_stq_idx(input rob_valids[63:0], input rob_uses_stq[63:0], input [3:0] rob_stq_indexes[63:0]);
	  integer i;
	  reg [15:0] stq_idx_used;
		begin
	    stq_idx_used = 16'b0;
	    for(i=0; i<=63; i=i+1)begin
	      if(rob_valids[i] && rob_uses_stq[i])
	      begin
		if(stq_idx_used[rob_stq_indexes[i]] == 1'b0)
		begin
		  stq_idx_used[rob_stq_indexes[i]] = 1'b1;
		end
		else
		begin
		  return 1'b0;
		end
	      end
	    end
	    return 1'b1;
		end
	endfunction
	
	wire unique_stq_idx_1;
	assign unique_stq_idx_1 = check_uniqueness_stq_idx(rob_valids_1, rob_uses_stq_1, rob_stq_indexes_1);*/
	
	wire stdf_clr_bsy_uses_stq_1;
	assign stdf_clr_bsy_uses_stq_1 = soc1.lsu.stdf_clr_bsy_valid ? rob_uses_stq_1[soc1.lsu.stdf_clr_bsy_rob_idx] : 1'b1;
	
	wire fdivsqrt_consistency_1;
	assign fdivsqrt_consistency_1 =
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val
	?
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A != 3'b0
	?
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B == 4'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C == 3'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E == 3'b0)
	:
	  1'b1
	) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B != 4'b0
	?
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A == 3'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C == 3'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E == 3'b0)
	:
	  1'b1
	) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C != 3'b0
	?
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B == 4'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A == 3'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E == 3'b0)
	:
	  1'b1
	) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E != 3'b0
	?
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B == 4'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C == 3'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A == 3'b0)
	:
	  1'b1
	) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PA
	?
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PB == 1'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PC == 1'b0)
	:
	  1'b1
	) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PB
	?
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PA == 1'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PC == 1'b0)
	:
	  1'b1
	) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PC
	?
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PB == 1'b0) &&
	  (soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PA == 1'b0)
	:
	  1'b1
	)
	:
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A == 3'b0) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B == 4'b0) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C == 3'b0) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E == 3'b0) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PA == 1'b0) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PB == 1'b0) &&
	(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PC == 1'b0)
	);
	
	wire unique_write_port_addr_1;
	assign unique_write_port_addr_1 =
		(soc1.core.iregfile.io_write_ports_0_valid && soc1.core.iregfile.io_write_ports_1_valid ? soc1.core.iregfile.io_write_ports_0_bits_addr != soc1.core.iregfile.io_write_ports_1_bits_addr : 1'b1) &&
		(soc1.core.iregfile.io_write_ports_0_valid && soc1.core.iregfile.io_write_ports_2_valid ? soc1.core.iregfile.io_write_ports_0_bits_addr != soc1.core.iregfile.io_write_ports_2_bits_addr : 1'b1) &&
		(soc1.core.iregfile.io_write_ports_1_valid && soc1.core.iregfile.io_write_ports_2_valid ? soc1.core.iregfile.io_write_ports_1_bits_addr != soc1.core.iregfile.io_write_ports_2_bits_addr : 1'b1)
	;
	
	wire lsu_req_consistent_1;
	assign lsu_req_consistent_1 =
		soc1.lsu.io_core_exe_0_req_valid
		?
			(soc1.lsu.io_core_exe_0_req_bits_uop_ctrl_is_load == soc1.lsu.io_core_exe_0_req_bits_uop_uses_ldq) &&
			((soc1.lsu.io_core_exe_0_req_bits_uop_ctrl_is_sta || soc1.lsu.io_core_exe_0_req_bits_uop_ctrl_is_std) == soc1.lsu.io_core_exe_0_req_bits_uop_uses_stq)
		:
			1'b1;
			
	wire csr_req_not_speculative_1;
	assign csr_req_not_speculative_1 = soc1.core.csr_exe_unit.io_req_valid && soc1.core.csr_exe_unit.io_req_bits_uop_ctrl_csr_cmd != 3'b0 ? soc1.core.csr_exe_unit.io_req_bits_uop_br_mask == 12'b0 : 1'b1;
	
	wire lsu_req_uses_queue_1;
	assign lsu_req_uses_queue_1 = soc1.lsu.io_core_exe_0_req_valid ? soc1.lsu.io_core_exe_0_req_bits_uop_uses_ldq || soc1.lsu.io_core_exe_0_req_bits_uop_uses_stq || (soc1.lsu.io_core_exe_0_req_bits_sfence_valid && soc1.lsu.io_core_exe_0_req_bits_uop_br_mask == 12'b0): 1'b1;
	
	wire dmem_resp_amo_1;
	assign dmem_resp_amo_1 =
	soc1.lsu.io_dmem_resp_0_valid && soc1.lsu.io_dmem_resp_0_bits_uop_is_amo
	?
		soc1.lsu.io_dmem_resp_0_bits_uop_uses_stq && stq_valids_1[soc1.lsu.io_dmem_resp_0_bits_uop_stq_idx] &&
		(rob_branch_masks_1[stq_rob_idx_1[soc1.lsu.io_dmem_resp_0_bits_uop_stq_idx]] == 12'b0) &&
		!stq_committed_1[soc1.lsu.io_dmem_resp_0_bits_uop_stq_idx] &&
		soc1.lsu.stq_head == soc1.lsu.io_dmem_resp_0_bits_uop_stq_idx &&
		soc1.core.rob.io_rob_head_idx == stq_rob_idx_1[soc1.lsu.io_dmem_resp_0_bits_uop_stq_idx] &&
		soc1.core.rob.io_rob_tail_idx == ((stq_rob_idx_1[soc1.lsu.io_dmem_resp_0_bits_uop_stq_idx] + 1) % 64)
	:
		1'b1
	;
	
	wire buffers_equal_STQ_1;
	assign buffers_equal_STQ_1 = 
		(soc1.lsu.fired_stdf_incoming && !stq_committed_1[soc1.lsu.mem_stdf_uop_stq_idx] ? stq_valids_1[soc1.lsu.mem_stdf_uop_stq_idx] && soc1.lsu.mem_stdf_uop_rob_idx == stq_rob_idx_1[soc1.lsu.mem_stdf_uop_stq_idx] : 1'b1) &&
		(soc1.core.iregister_read.exe_reg_valids_0 && soc1.core.iregister_read.exe_reg_uops_0_uses_stq && !stq_committed_1[soc1.core.iregister_read.exe_reg_uops_0_stq_idx] ? stq_valids_1[soc1.core.iregister_read.exe_reg_uops_0_stq_idx] && soc1.core.iregister_read.exe_reg_uops_0_rob_idx == stq_rob_idx_1[soc1.core.iregister_read.exe_reg_uops_0_stq_idx] : 1'b1);
	
	wire buffers_equal_LDQ_1;
	assign buffers_equal_LDQ_1 =
	  (soc1.core.iregister_read.exe_reg_valids_0 && soc1.core.iregister_read.exe_reg_uops_0_uses_ldq ? ldq_valids_1[soc1.core.iregister_read.exe_reg_uops_0_ldq_idx] && soc1.core.iregister_read.exe_reg_uops_0_rob_idx == ldq_rob_idx_1[soc1.core.iregister_read.exe_reg_uops_0_ldq_idx] : 1'b1);

	
	wire ldq_head_empty_1;
	assign ldq_head_empty_1 = !ldq_valids_1[soc1.lsu.ldq_head] == (!ldq_valids_1[0] && !ldq_valids_1[1] && !ldq_valids_1[2] && !ldq_valids_1[3] && !ldq_valids_1[4] && !ldq_valids_1[5] && !ldq_valids_1[6] && !ldq_valids_1[7] && !ldq_valids_1[8] &&
	 !ldq_valids_1[9] && !ldq_valids_1[10] && !ldq_valids_1[11] && !ldq_valids_1[12] && !ldq_valids_1[13] && !ldq_valids_1[14] && !ldq_valids_1[15]);


	function automatic check_uniqueness_ldq_rob_idx(input ldq_valids[15:0], input [5:0] ldq_rob_idx[15:0]);
	  integer i;
	  reg [63:0] rob_idx_used;
	  begin
	    rob_idx_used = 64'b0;
	    for(i=0; i<=15; i=i+1)begin
	      if(ldq_valids[i])
	      begin
	  if(rob_idx_used[ldq_rob_idx[i]] == 1'b0)
	  begin
	    rob_idx_used[ldq_rob_idx[i]] = 1'b1;
	  end
	  else
	  begin
	    return 1'b0;
	  end
	      end
	    end
	    return 1'b1;
	  end
	endfunction
	
	wire unique_ldq_rob_idx_1;
	assign unique_ldq_rob_idx_1 = check_uniqueness_ldq_rob_idx(ldq_valids_1, ldq_rob_idx_1);
	
	/*wire mem_xcpt_consistency_1;
	assign mem_xcpt_consistency_1 =
	  soc1.lsu.will_fire_store_commit_0 && soc1.lsu.mem_xcpt_valids_0
	  ?
	    soc1.lsu.mem_xcpt_uops_0_stq_idx == soc1.lsu.stq_execute_head && soc1.lsu.mem_xcpt_uops_0_uses_stq
	  :
	    1'b1;*/
	
	wire fired_load_incoming_conflicts_1;
	assign fired_load_incoming_conflicts_1 =
	  !(soc1.lsu.fired_load_incoming_REG && soc1.lsu.fired_stad_incoming_REG) &&
	  !(soc1.lsu.fired_load_incoming_REG && soc1.lsu.fired_sta_incoming_REG) &&
	  !(soc1.lsu.fired_load_incoming_REG && soc1.lsu.fired_sfence_0) &&
	  !(soc1.lsu.fired_load_incoming_REG && soc1.lsu.fired_load_retry_REG) &&
	  !(soc1.lsu.fired_load_incoming_REG && soc1.lsu.fired_sta_retry_REG) &&
	  !(soc1.lsu.fired_load_incoming_REG && soc1.lsu.fired_release_0) &&
	  !(soc1.lsu.fired_load_incoming_REG && soc1.lsu.fired_load_wakeup_REG);
	  
	wire fired_stad_incoming_conflicts_1;
	assign fired_stad_incoming_conflicts_1 =
	  !(soc1.lsu.fired_stad_incoming_REG && soc1.lsu.fired_sta_incoming_REG) &&
	  !(soc1.lsu.fired_stad_incoming_REG && soc1.lsu.fired_std_incoming_REG) &&
	  !(soc1.lsu.fired_stad_incoming_REG && soc1.lsu.fired_sfence_0) &&
	  !(soc1.lsu.fired_stad_incoming_REG && soc1.lsu.fired_release_0) &&
	  !(soc1.lsu.fired_stad_incoming_REG && soc1.lsu.fired_load_retry_REG) &&
	  !(soc1.lsu.fired_stad_incoming_REG && soc1.lsu.fired_sta_retry_REG) &&
	  !(soc1.lsu.fired_stad_incoming_REG && soc1.lsu.fired_load_wakeup_REG);

	wire fired_sta_incoming_conflicts_1;
	assign fired_sta_incoming_conflicts_1 =
	  !(soc1.lsu.fired_sta_incoming_REG && soc1.lsu.fired_std_incoming_REG) &&
	  !(soc1.lsu.fired_sta_incoming_REG && soc1.lsu.fired_sfence_0) &&
	  !(soc1.lsu.fired_sta_incoming_REG && soc1.lsu.fired_release_0) &&
	  !(soc1.lsu.fired_sta_incoming_REG && soc1.lsu.fired_load_retry_REG) &&
	  !(soc1.lsu.fired_sta_incoming_REG && soc1.lsu.fired_sta_retry_REG) &&
	  !(soc1.lsu.fired_sta_incoming_REG && soc1.lsu.fired_load_wakeup_REG);

	wire fired_std_incoming_conflicts_1;
	assign fired_std_incoming_conflicts_1 =
	  !(soc1.lsu.fired_std_incoming_REG && soc1.lsu.fired_sfence_0) &&
	  !(soc1.lsu.fired_std_incoming_REG && soc1.lsu.fired_sta_retry_REG);

	wire fired_std_conflicts_1;
	assign fired_std_conflicts_1 =
	  1'b1;

	wire fired_sfence_conflicts_1;
	assign fired_sfence_conflicts_1 = 
	  !(soc1.lsu.fired_sfence_0 && soc1.lsu.fired_load_retry_REG) &&
	  !(soc1.lsu.fired_sfence_0 && soc1.lsu.fired_sta_retry_REG);

	wire fired_release_conflicts_1;
	assign fired_release_conflicts_1 = 
	  !(soc1.lsu.fired_release_0 && soc1.lsu.fired_load_retry_REG) &&
	  !(soc1.lsu.fired_release_0 && soc1.lsu.fired_sta_retry_REG);

	wire fired_load_retry_conflicts_1;
	assign fired_load_retry_conflicts_1 = 
	  !(soc1.lsu.fired_load_retry_REG && soc1.lsu.fired_sta_retry_REG) &&
	  !(soc1.lsu.fired_load_retry_REG && soc1.lsu.fired_load_wakeup_REG);

	wire fired_sta_retry_conflicts_1;
	assign fired_sta_retry_conflicts_1 = 
	  !(soc1.lsu.fired_sta_retry_REG && soc1.lsu.fired_load_wakeup_REG);
	
	function automatic check_uopc_lrs1_lrs2(input [6:0] uopc, input [1:0] lrs1_type, input [1:0] lrs2_type);
	begin
	  case (uopc)
	  7'h0 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopNOP
	  7'h1 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopLD
	  7'h2 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2 || lrs2_type == 2'h0); // uopSTA
	  7'h3 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h0); // uopSTD
	  7'h4 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopLUI
	  7'h5 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopADDI
	  7'h6 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopANDI
	  7'h7 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopORI
	  7'h8 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopXORI
	  7'h9 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSLTI
	  7'ha : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSLTIU
	  7'hb : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSLLI
	  7'hc : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRAI
	  7'hd : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRLI
	  7'he : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSLL
	  7'hf : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopADD
	  7'h10 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSUB
	  7'h11 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSLT
	  7'h12 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSLTU
	  7'h13 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopAND
	  7'h14 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopOR
	  7'h15 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopXOR
	  7'h16 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSRA
	  7'h17 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSRL
	  7'h18 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBEQ
	  7'h19 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBNE
	  7'h1a : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBGE
	  7'h1b : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBGEU
	  7'h1c : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBLT
	  7'h1d : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBLTU
	  7'h1e : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopCSRRW
	  7'h1f : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopCSRRS
	  7'h20 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopCSRRC
	  7'h21 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h3) && (lrs2_type == 2'h2); // uopCSRRWI
	  7'h22 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h3) && (lrs2_type == 2'h2); // uopCSRRSI
	  7'h23 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h3) && (lrs2_type == 2'h2); // uopCSRRCI
	  //7'h24 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopJ
	  7'h25 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopJAL
	  7'h26 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopJALR
	  7'h27 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopAUIPC
	  //7'h28 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRET
	  //7'h29 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopCFLSH
	  7'h2a : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopFENCE
	  7'h2b : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopADDIW
	  7'h2c : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopADDW
	  7'h2d : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSUBW
	  7'h2e : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSLLIW
	  7'h2f : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSLLW
	  7'h30 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRAIW
	  7'h31 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSRAW
	  7'h32 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRLIW
	  7'h33 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSRLW
	  7'h34 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMUL
	  7'h35 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMULH
	  7'h36 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMULHU
	  7'h37 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMULHSU
	  7'h38 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMULW
	  7'h39 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopDIV
	  7'h3a : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopDIVU
	  7'h3b : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopREM
	  7'h3c : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopREMU
	  7'h3d : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopDIVW
	  7'h3e : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopDIVUW
	  7'h3f : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopREMW
	  7'h40 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopREMUW
	  //7'h41 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFENCEI
	  //7'h42 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // XXXXXXXXX
	  7'h43 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopAMO_AG
	  7'h44 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFMV_S_X
	  7'h45 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFMV_D_X
	  7'h46 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFMV_X_S
	  7'h47 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFMV_X_D
	  7'h48 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFSGNJ_S
	  7'h49 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFSGNJ_D
	  7'h4a : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCVT_S_D
	  7'h4b : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCVT_D_S
	  7'h4c : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFCVT_S_X
	  7'h4d : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFCVT_D_X
	  7'h4e : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCVT_X_S
	  7'h4f : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCVT_X_D
	  7'h50 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopCMPR_S
	  7'h51 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopCMPR_D
	  7'h52 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCLASS_S
	  7'h53 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCLASS_D
	  7'h54 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMINMAX_S
	  7'h55 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMINMAX_D
	  //7'h56 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // XXXXXXXXX
	  7'h57 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFADD_S
	  7'h58 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFSUB_S
	  7'h59 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMUL_S
	  7'h5a : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFADD_D
	  7'h5b : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFSUB_D
	  7'h5c : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMUL_D
	  7'h5d : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMADD_S
	  7'h5e : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMSUB_S
	  7'h5f : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFNMADD_S
	  7'h60 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFNMSUB_S
	  7'h61 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMADD_D
	  7'h62 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMSUB_D
	  7'h63 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFNMADD_D
	  7'h64 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFNMSUB_D
	  7'h65 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFDIV_S
	  7'h66 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFDIV_D
	  7'h67 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFSQRT_S
	  7'h68 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFSQRT_D
	  7'h69 : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopWFI
	  7'h6a : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopERET
	  7'h6b : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSFENCE
	  7'h6c : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0 || lrs1_type == 2'h2) && (lrs2_type == 2'h0 || lrs2_type == 2'h2); // uopROCC
	  //7'h6d : check_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopMOV
	   default : check_uopc_lrs1_lrs2 = 1'b0;
	  endcase
	end
	endfunction

	function automatic check_fp_uopc_lrs1_lrs2(input [6:0] uopc, input [1:0] lrs1_type, input [1:0] lrs2_type);
	begin
	  case (uopc)
	  7'h0 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopNOP
	  7'h1 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopLD
	  7'h2 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h1); // uopSTA
	  7'h3 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h0); // uopSTD
	  7'h4 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopLUI
	  7'h5 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopADDI
	  7'h6 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopANDI
	  7'h7 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopORI
	  7'h8 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopXORI
	  7'h9 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSLTI
	  7'ha : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSLTIU
	  7'hb : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSLLI
	  7'hc : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRAI
	  7'hd : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRLI
	  7'he : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSLL
	  7'hf : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopADD
	  7'h10 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSUB
	  7'h11 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSLT
	  7'h12 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSLTU
	  7'h13 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopAND
	  7'h14 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopOR
	  7'h15 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopXOR
	  7'h16 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSRA
	  7'h17 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSRL
	  7'h18 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBEQ
	  7'h19 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBNE
	  7'h1a : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBGE
	  7'h1b : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBGEU
	  7'h1c : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBLT
	  7'h1d : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopBLTU
	  7'h1e : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopCSRRW
	  7'h1f : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopCSRRS
	  7'h20 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopCSRRC
	  7'h21 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h3) && (lrs2_type == 2'h2); // uopCSRRWI
	  7'h22 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h3) && (lrs2_type == 2'h2); // uopCSRRSI
	  7'h23 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h3) && (lrs2_type == 2'h2); // uopCSRRCI
	  //7'h24 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopJ
	  7'h25 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopJAL
	  7'h26 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopJALR
	  7'h27 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopAUIPC
	  //7'h28 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRET
	  //7'h29 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopCFLSH
	  7'h2a : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopFENCE
	  7'h2b : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopADDIW
	  7'h2c : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopADDW
	  7'h2d : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSUBW
	  7'h2e : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSLLIW
	  7'h2f : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSLLW
	  7'h30 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRAIW
	  7'h31 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSRAW
	  7'h32 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopSRLIW
	  7'h33 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSRLW
	  7'h34 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMUL
	  7'h35 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMULH
	  7'h36 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMULHU
	  7'h37 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMULHSU
	  7'h38 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopMULW
	  7'h39 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopDIV
	  7'h3a : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopDIVU
	  7'h3b : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopREM
	  7'h3c : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopREMU
	  7'h3d : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopDIVW
	  7'h3e : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopDIVUW
	  7'h3f : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopREMW
	  7'h40 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopREMUW
	  //7'h41 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFENCEI
	  //7'h42 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // XXXXXXXXX
	  7'h43 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopAMO_AG
	  7'h44 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFMV_S_X
	  7'h45 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFMV_D_X
	  7'h46 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFMV_X_S
	  7'h47 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFMV_X_D
	  7'h48 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFSGNJ_S
	  7'h49 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFSGNJ_D
	  7'h4a : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCVT_S_D
	  7'h4b : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCVT_D_S
	  7'h4c : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFCVT_S_X
	  7'h4d : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopFCVT_D_X
	  7'h4e : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCVT_X_S
	  7'h4f : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCVT_X_D
	  7'h50 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopCMPR_S
	  7'h51 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopCMPR_D
	  7'h52 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCLASS_S
	  7'h53 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFCLASS_D
	  7'h54 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMINMAX_S
	  7'h55 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMINMAX_D
	  //7'h56 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // XXXXXXXXX
	  7'h57 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFADD_S
	  7'h58 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFSUB_S
	  7'h59 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMUL_S
	  7'h5a : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFADD_D
	  7'h5b : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFSUB_D
	  7'h5c : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMUL_D
	  7'h5d : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMADD_S
	  7'h5e : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMSUB_S
	  7'h5f : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFNMADD_S
	  7'h60 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFNMSUB_S
	  7'h61 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMADD_D
	  7'h62 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFMSUB_D
	  7'h63 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFNMADD_D
	  7'h64 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFNMSUB_D
	  7'h65 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFDIV_S
	  7'h66 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h1); // uopFDIV_D
	  7'h67 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFSQRT_S
	  7'h68 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h1) && (lrs2_type == 2'h2); // uopFSQRT_D
	  7'h69 : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopWFI
	  7'h6a : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h2) && (lrs2_type == 2'h2); // uopERET
	  7'h6b : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h0); // uopSFENCE
	  7'h6c : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0 || lrs1_type == 2'h2) && (lrs2_type == 2'h0 || lrs2_type == 2'h2); // uopROCC
	  //7'h6d : check_fp_uopc_lrs1_lrs2 = (lrs1_type == 2'h0) && (lrs2_type == 2'h2); // uopMOV
	   default : check_fp_uopc_lrs1_lrs2 = 1'b0;
	  endcase
	end
	endfunction
	    
	wire rrd_lrs_types_1;
	assign rrd_lrs_types_1 =
	check_uopc_lrs1_lrs2(soc1.core.iregister_read.rrd_uops_0_REG_uopc, soc1.core.iregister_read.rrd_uops_0_REG_lrs1_rtype, soc1.core.iregister_read.rrd_uops_0_REG_lrs2_rtype) &&
	check_uopc_lrs1_lrs2(soc1.core.iregister_read.rrd_uops_1_REG_uopc, soc1.core.iregister_read.rrd_uops_1_REG_lrs1_rtype, soc1.core.iregister_read.rrd_uops_1_REG_lrs2_rtype) &&
	check_uopc_lrs1_lrs2(soc1.core.iregister_read.rrd_uops_2_REG_uopc, soc1.core.iregister_read.rrd_uops_2_REG_lrs1_rtype, soc1.core.iregister_read.rrd_uops_2_REG_lrs2_rtype) &&
	check_fp_uopc_lrs1_lrs2(soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uopc, soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_lrs1_rtype, soc1.core.fp_pipeline.fregister_read.rrd_uops_0_REG_lrs2_rtype);
	
	
	function automatic check_uopc_op_sel(input [6:0] uopc, input [1:0] op1_sel, input [2:0] op2_sel);
	begin
	  case (uopc)
	  7'h0 : check_uopc_op_sel = 1'b1; // uopNOP
	  7'h1 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopLD
	  7'h2 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopSTA
	  7'h3 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSTD
	  7'h4 : check_uopc_op_sel = (op1_sel == 2'h1) && (op2_sel == 3'h1); // uopLUI
	  7'h5 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopADDI
	  7'h6 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopANDI
	  7'h7 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopORI
	  7'h8 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopXORI
	  7'h9 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopSLTI
	  7'ha : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopSLTIU
	  7'hb : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopSLLI
	  7'hc : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopSRAI
	  7'hd : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopSRLI
	  7'he : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSLL
	  7'hf : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopADD
	  7'h10 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSUB
	  7'h11 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSLT
	  7'h12 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSLTU
	  7'h13 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopAND
	  7'h14 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopOR
	  7'h15 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopXOR
	  7'h16 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSRA
	  7'h17 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSRL
	  7'h18 : check_uopc_op_sel = 1'b1; // uopBEQ
	  7'h19 : check_uopc_op_sel = 1'b1; // uopBNE
	  7'h1a : check_uopc_op_sel = 1'b1; // uopBGE
	  7'h1b : check_uopc_op_sel = 1'b1; // uopBGEU
	  7'h1c : check_uopc_op_sel = 1'b1; // uopBLT
	  7'h1d : check_uopc_op_sel = 1'b1; // uopBLTU
	  7'h1e : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h2); // uopCSRRW
	  7'h1f : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h2); // uopCSRRS
	  7'h20 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h2); // uopCSRRC
	  7'h21 : check_uopc_op_sel = (op1_sel == 2'h1) && (op2_sel == 3'h4); // uopCSRRWI
	  7'h22 : check_uopc_op_sel = (op1_sel == 2'h1) && (op2_sel == 3'h4); // uopCSRRSI
	  7'h23 : check_uopc_op_sel = (op1_sel == 2'h1) && (op2_sel == 3'h4); // uopCSRRCI
	  //7'h24 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 2'h2); // uopJ
	  7'h25 : check_uopc_op_sel = (op1_sel == 2'h2) && (op2_sel == 3'h3); // uopJAL
	  7'h26 : check_uopc_op_sel = (op1_sel == 2'h2) && (op2_sel == 3'h3); // uopJALR
	  7'h27 : check_uopc_op_sel = (op1_sel == 2'h2) && (op2_sel == 3'h1); // uopAUIPC
	  //7'h28 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 2'h2); // uopSRET
	  //7'h29 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 2'h2); // uopCFLSH
	  7'h2a : check_uopc_op_sel = 1'b1; // uopFENCE
	  7'h2b : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopADDIW
	  7'h2c : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopADDW
	  7'h2d : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSUBW
	  7'h2e : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopSLLIW
	  7'h2f : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSLLW
	  7'h30 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopSRAIW
	  7'h31 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSRAW
	  7'h32 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h1); // uopSRLIW
	  7'h33 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSRLW
	  7'h34 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopMUL
	  7'h35 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopMULH
	  7'h36 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopMULHU
	  7'h37 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopMULHSU
	  7'h38 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopMULW
	  7'h39 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopDIV
	  7'h3a : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopDIVU
	  7'h3b : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopREM
	  7'h3c : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopREMU
	  7'h3d : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopDIVW
	  7'h3e : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopDIVUW
	  7'h3f : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopREMW
	  7'h40 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopREMUW
	  //7'h41 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 2'h2); // uopFENCEI
	  //7'h42 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 2'h2); // XXXXXXXXX
	  7'h43 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h2); // uopAMO_AG
	  7'h44 : check_uopc_op_sel = 1'b1; // uopFMV_S_X
	  7'h45 : check_uopc_op_sel = 1'b1; // uopFMV_D_X
	  7'h46 : check_uopc_op_sel = 1'b1; // uopFMV_X_S
	  7'h47 : check_uopc_op_sel = 1'b1; // uopFMV_X_D
	  7'h48 : check_uopc_op_sel = 1'b1; // uopFSGNJ_S
	  7'h49 : check_uopc_op_sel = 1'b1; // uopFSGNJ_D
	  7'h4a : check_uopc_op_sel = 1'b1; // uopFCVT_S_D
	  7'h4b : check_uopc_op_sel = 1'b1; // uopFCVT_D_S
	  7'h4c : check_uopc_op_sel = 1'b1; // uopFCVT_S_X
	  7'h4d : check_uopc_op_sel = 1'b1; // uopFCVT_D_X
	  7'h4e : check_uopc_op_sel = 1'b1; // uopFCVT_X_S
	  7'h4f : check_uopc_op_sel = 1'b1; // uopFCVT_X_D
	  7'h50 : check_uopc_op_sel = 1'b1; // uopCMPR_S
	  7'h51 : check_uopc_op_sel = 1'b1; // uopCMPR_D
	  7'h52 : check_uopc_op_sel = 1'b1; // uopFCLASS_S
	  7'h53 : check_uopc_op_sel = 1'b1; // uopFCLASS_D
	  7'h54 : check_uopc_op_sel = 1'b1; // uopFMINMAX_S
	  7'h55 : check_uopc_op_sel = 1'b1; // uopFMINMAX_D
	  //7'h56 : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 2'h2); // XXXXXXXXX
	  7'h57 : check_uopc_op_sel = 1'b1; // uopFADD_S
	  7'h58 : check_uopc_op_sel = 1'b1; // uopFSUB_S
	  7'h59 : check_uopc_op_sel = 1'b1; // uopFMUL_S
	  7'h5a : check_uopc_op_sel = 1'b1; // uopFADD_D
	  7'h5b : check_uopc_op_sel = 1'b1; // uopFSUB_D
	  7'h5c : check_uopc_op_sel = 1'b1; // uopFMUL_D
	  7'h5d : check_uopc_op_sel = 1'b1; // uopFMADD_S
	  7'h5e : check_uopc_op_sel = 1'b1; // uopFMSUB_S
	  7'h5f : check_uopc_op_sel = 1'b1; // uopFNMADD_S
	  7'h60 : check_uopc_op_sel = 1'b1; // uopFNMSUB_S
	  7'h61 : check_uopc_op_sel = 1'b1; // uopFMADD_D
	  7'h62 : check_uopc_op_sel = 1'b1; // uopFMSUB_D
	  7'h63 : check_uopc_op_sel = 1'b1; // uopFNMADD_D
	  7'h64 : check_uopc_op_sel = 1'b1; // uopFNMSUB_D
	  7'h65 : check_uopc_op_sel = 1'b1; // uopFDIV_S
	  7'h66 : check_uopc_op_sel = 1'b1; // uopFDIV_D
	  7'h67 : check_uopc_op_sel = 1'b1; // uopFSQRT_S
	  7'h68 : check_uopc_op_sel = 1'b1; // uopFSQRT_D
	  7'h69 : check_uopc_op_sel = (op1_sel == 2'h1) && (op2_sel == 3'h4); // uopWFI
	  7'h6a : check_uopc_op_sel = (op1_sel == 2'h1) && (op2_sel == 3'h4); // uopERET
	  7'h6b : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 3'h0); // uopSFENCE
	  7'h6c : check_uopc_op_sel = 1'b1; // uopROCC
	  //7'h6d : check_uopc_op_sel = (op1_sel == 2'h0) && (op2_sel == 2'h2); // uopMOV
	   default : check_uopc_op_sel = 1'b0;
	  endcase
	end
	endfunction
	
	wire rrd_op_sel_1;
	assign rrd_op_sel_1 =
		check_uopc_op_sel(soc1.core.iregister_read.rrd_uops_1_REG_uopc, soc1.core.iregister_read.rrd_uops_1_REG_ctrl_op1_sel, soc1.core.iregister_read.rrd_uops_1_REG_ctrl_op2_sel) &&
		check_uopc_op_sel(soc1.core.iregister_read.rrd_uops_2_REG_uopc, soc1.core.iregister_read.rrd_uops_2_REG_ctrl_op1_sel, soc1.core.iregister_read.rrd_uops_2_REG_ctrl_op2_sel);
	
	function automatic check_csr_alu_uopc(input [6:0] uopc);
	begin
	  case (uopc)
	    7'hb  : check_csr_alu_uopc = 1'b1; // uopSLLI
	    7'hd  : check_csr_alu_uopc = 1'b1; // uopSRLI
	    7'hc  : check_csr_alu_uopc = 1'b1; // uopSRAI
	    7'h2b : check_csr_alu_uopc = 1'b1; // uopADDIW
	    7'h2e : check_csr_alu_uopc = 1'b1; // uopSLLIW
	    7'h30 : check_csr_alu_uopc = 1'b1; // uopSRAIW
	    7'h32 : check_csr_alu_uopc = 1'b1; // uopSRLIW
	    7'h2c : check_csr_alu_uopc = 1'b1; // uopADDW
	    7'h2d : check_csr_alu_uopc = 1'b1; // uopSUBW
	    7'h2f : check_csr_alu_uopc = 1'b1; // uopSLLW
	    7'h31 : check_csr_alu_uopc = 1'b1; // uopSRAW
	    7'h33 : check_csr_alu_uopc = 1'b1; // uopSRLW
	    7'h4  : check_csr_alu_uopc = 1'b1; // uopLUI
	    7'h5  : check_csr_alu_uopc = 1'b1; // uopADDI
	    7'h6  : check_csr_alu_uopc = 1'b1; // uopANDI
	    7'h7  : check_csr_alu_uopc = 1'b1; // uopORI
	    7'h8  : check_csr_alu_uopc = 1'b1; // uopXORI
	    7'h9  : check_csr_alu_uopc = 1'b1; // uopSLTI
	    7'ha  : check_csr_alu_uopc = 1'b1; // uopSLTIU
	    7'he  : check_csr_alu_uopc = 1'b1; // uopSLL
	    7'hf  : check_csr_alu_uopc = 1'b1; // uopADD
	    7'h10 : check_csr_alu_uopc = 1'b1; // uopSUB
	    7'h11 : check_csr_alu_uopc = 1'b1; // uopSLT
	    7'h12 : check_csr_alu_uopc = 1'b1; // uopSLTU
	    7'h13 : check_csr_alu_uopc = 1'b1; // uopAND
	    7'h14 : check_csr_alu_uopc = 1'b1; // uopOR
	    7'h15 : check_csr_alu_uopc = 1'b1; // uopXOR
	    7'h16 : check_csr_alu_uopc = 1'b1; // uopSRA
	    7'h17 : check_csr_alu_uopc = 1'b1; // uopSRL
	    7'h18 : check_csr_alu_uopc = 1'b1; // uopBEQ
	    7'h19 : check_csr_alu_uopc = 1'b1; // uopBNE
	    7'h1a : check_csr_alu_uopc = 1'b1; // uopBGE
	    7'h1b : check_csr_alu_uopc = 1'b1; // uopBGEU
	    7'h1c : check_csr_alu_uopc = 1'b1; // uopBLT
	    7'h1d : check_csr_alu_uopc = 1'b1; // uopBLTU
	    7'h27 : check_csr_alu_uopc = 1'b1; // uopAUIPC
	    7'h25 : check_csr_alu_uopc = 1'b1; // uopJAL
	    7'h26 : check_csr_alu_uopc = 1'b1; // uopJALR
	    7'h1e : check_csr_alu_uopc = 1'b1; // uopCSRRW
	    7'h1f : check_csr_alu_uopc = 1'b1; // uopCSRRS
	    7'h20 : check_csr_alu_uopc = 1'b1; // uopCSRRC
	    7'h21 : check_csr_alu_uopc = 1'b1; // uopCSRRWI
	    7'h22 : check_csr_alu_uopc = 1'b1; // uopCSRRSI
	    7'h23 : check_csr_alu_uopc = 1'b1; // uopCSRRCI
	    7'h6a : check_csr_alu_uopc = 1'b1; // uopERET
	    7'h69 : check_csr_alu_uopc = 1'b1; // uopWFI
	    7'h6c : check_csr_alu_uopc = 1'b1; // uopROCC
	    default : check_csr_alu_uopc = 1'b0;
	  endcase
	end
	endfunction
	
	wire csr_alu_req_uopc_1;
	assign csr_alu_req_uopc_1 = !soc1.core.csr_exe_unit.alu.io_req_valid || check_csr_alu_uopc(soc1.core.csr_exe_unit.alu.io_req_bits_uop_uopc);
	
	function automatic check_csr_div_uopc(input [6:0] uopc);
	begin
	  case (uopc)
	    7'h39 : check_csr_div_uopc = 1'b1; // uopDIV
	    7'h3a : check_csr_div_uopc = 1'b1; // uopDIVU
	    7'h3b : check_csr_div_uopc = 1'b1; // uopREM
	    7'h3c : check_csr_div_uopc = 1'b1; // uopREMU
	    7'h3d : check_csr_div_uopc = 1'b1; // uopDIVW
	    7'h3e : check_csr_div_uopc = 1'b1; // uopDIVUW
	    7'h3f : check_csr_div_uopc = 1'b1; // uopREMW
	    7'h40 : check_csr_div_uopc = 1'b1; // uopREMUW
	    default : check_csr_div_uopc = 1'b0;
	  endcase
	end
	endfunction
	
	wire csr_div_req_uopc_1;
	assign csr_div_req_uopc_1 = !soc1.core.csr_exe_unit.div.io_req_valid || check_csr_div_uopc(soc1.core.csr_exe_unit.div.io_req_bits_uop_uopc);
	
	function automatic check_jmp_unit_alu_uopc(input [6:0] uopc);
	begin
	  case (uopc)
	    7'hb  : check_jmp_unit_alu_uopc = 1'b1; // uopSLLI
	    7'hd  : check_jmp_unit_alu_uopc = 1'b1; // uopSRLI
	    7'hc  : check_jmp_unit_alu_uopc = 1'b1; // uopSRAI
	    7'h2b : check_jmp_unit_alu_uopc = 1'b1; // uopADDIW
	    7'h2e : check_jmp_unit_alu_uopc = 1'b1; // uopSLLIW
	    7'h30 : check_jmp_unit_alu_uopc = 1'b1; // uopSRAIW
	    7'h32 : check_jmp_unit_alu_uopc = 1'b1; // uopSRLIW
	    7'h2c : check_jmp_unit_alu_uopc = 1'b1; // uopADDW
	    7'h2d : check_jmp_unit_alu_uopc = 1'b1; // uopSUBW
	    7'h2f : check_jmp_unit_alu_uopc = 1'b1; // uopSLLW
	    7'h31 : check_jmp_unit_alu_uopc = 1'b1; // uopSRAW
	    7'h33 : check_jmp_unit_alu_uopc = 1'b1; // uopSRLW
	    7'h4  : check_jmp_unit_alu_uopc = 1'b1; // uopLUI
	    7'h5  : check_jmp_unit_alu_uopc = 1'b1; // uopADDI
	    7'h6  : check_jmp_unit_alu_uopc = 1'b1; // uopANDI
	    7'h7  : check_jmp_unit_alu_uopc = 1'b1; // uopORI
	    7'h8  : check_jmp_unit_alu_uopc = 1'b1; // uopXORI
	    7'h9  : check_jmp_unit_alu_uopc = 1'b1; // uopSLTI
	    7'ha  : check_jmp_unit_alu_uopc = 1'b1; // uopSLTIU
	    7'he  : check_jmp_unit_alu_uopc = 1'b1; // uopSLL
	    7'hf  : check_jmp_unit_alu_uopc = 1'b1; // uopADD
	    7'h10 : check_jmp_unit_alu_uopc = 1'b1; // uopSUB
	    7'h11 : check_jmp_unit_alu_uopc = 1'b1; // uopSLT
	    7'h12 : check_jmp_unit_alu_uopc = 1'b1; // uopSLTU
	    7'h13 : check_jmp_unit_alu_uopc = 1'b1; // uopAND
	    7'h14 : check_jmp_unit_alu_uopc = 1'b1; // uopOR
	    7'h15 : check_jmp_unit_alu_uopc = 1'b1; // uopXOR
	    7'h16 : check_jmp_unit_alu_uopc = 1'b1; // uopSRA
	    7'h17 : check_jmp_unit_alu_uopc = 1'b1; // uopSRL
	    7'h18 : check_jmp_unit_alu_uopc = 1'b1; // uopBEQ
	    7'h19 : check_jmp_unit_alu_uopc = 1'b1; // uopBNE
	    7'h1a : check_jmp_unit_alu_uopc = 1'b1; // uopBGE
	    7'h1b : check_jmp_unit_alu_uopc = 1'b1; // uopBGEU
	    7'h1c : check_jmp_unit_alu_uopc = 1'b1; // uopBLT
	    7'h1d : check_jmp_unit_alu_uopc = 1'b1; // uopBLTU
	    7'h27 : check_jmp_unit_alu_uopc = 1'b1; // uopAUIPC
	    7'h25 : check_jmp_unit_alu_uopc = 1'b1; // uopJAL
	    7'h26 : check_jmp_unit_alu_uopc = 1'b1; // uopJALR
	    7'h1e : check_jmp_unit_alu_uopc = 1'b1; // uopCSRRW
	    7'h1f : check_jmp_unit_alu_uopc = 1'b1; // uopCSRRS
	    7'h20 : check_jmp_unit_alu_uopc = 1'b1; // uopCSRRC
	    7'h21 : check_jmp_unit_alu_uopc = 1'b1; // uopCSRRWI
	    7'h22 : check_jmp_unit_alu_uopc = 1'b1; // uopCSRRSI
	    7'h23 : check_jmp_unit_alu_uopc = 1'b1; // uopCSRRCI
	    7'h6a : check_jmp_unit_alu_uopc = 1'b1; // uopERET
	    7'h69 : check_jmp_unit_alu_uopc = 1'b1; // uopWFI
	    7'h6c : check_jmp_unit_alu_uopc = 1'b1; // uopROCC
	    default : check_jmp_unit_alu_uopc = 1'b0;
	  endcase
	end
	endfunction
	
	wire jmp_unit_alu_req_uopc_1;
	assign jmp_unit_alu_req_uopc_1 = !soc1.core.jmp_unit.alu.io_req_valid || check_jmp_unit_alu_uopc(soc1.core.jmp_unit.alu.io_req_bits_uop_uopc);
	
	wire dmem_resp_equals_s2_type_1;
	assign dmem_resp_equals_s2_type_1 = soc1.lsu.io_dmem_resp_0_valid && soc1.dcache.cache_resp_0_valid ? soc1.dcache.s2_type == 3'h4 || soc1.dcache.s2_type == 3'h0 : 1'b1;
	
	wire s2_hella_matching_s2_type_1;
	assign s2_hella_matching_s2_type_1 = soc1.dcache.s2_valid_REG && soc1.dcache.s2_req_0_is_hella ? soc1.dcache.s2_type == 3'h4 : 1'b1; 
	
	wire will_fire_sfence_not_speculative_1;
	assign will_fire_sfence_not_speculative_1 = soc1.lsu.will_fire_sfence_0_will_fire ? soc1.lsu.io_core_exe_0_req_bits_uop_br_mask == 12'h0 : 1'b1;

	wire store_req_not_committed_1;
	assign store_req_not_committed_1 = soc1.lsu.io_core_exe_0_req_valid && soc1.lsu.io_core_exe_0_req_bits_uop_uses_stq ? !stq_committed_1[soc1.lsu.io_core_exe_0_req_bits_uop_stq_idx] : 1'b1;
	
	wire hella_not_using_ldq_stq_1;
	assign hella_not_using_ldq_stq_1 = soc1.lsu.io_dmem_resp_0_bits_is_hella ? !soc1.lsu.io_dmem_resp_0_bits_uop_uses_ldq && !soc1.lsu.io_dmem_resp_0_bits_uop_uses_stq : 1'b1;
	
	wire s2_amo_nonspeculative_1;
	assign s2_amo_nonspeculative_1 = soc1.dcache.s2_valid_REG && soc1.dcache.s2_req_0_uop_is_amo ? soc1.dcache.s2_req_0_uop_br_mask == 12'h0 : 1'b1;
	
	wire committed_store_not_being_tainted_1;
	assign committed_store_not_being_tainted_1 =
		//GEN signals can be found by searching for io_core_exe_0_req_valid & io_core_exe_0_req_bits_uop_uses_stq & io_core_exe_0_req_bits_uop_taint ? _GEN_37623 : _GEN_37485; // @[lsu.scala 1580:89]
		(stq_valids_1[0] && stq_committed_1[0] ? !soc1.lsu._GEN_37477 : 1'b1) &&
		(stq_valids_1[1] && stq_committed_1[1] ? !soc1.lsu._GEN_37478 : 1'b1) &&
		(stq_valids_1[2] && stq_committed_1[2] ? !soc1.lsu._GEN_37479 : 1'b1) &&
		(stq_valids_1[3] && stq_committed_1[3] ? !soc1.lsu._GEN_37480 : 1'b1) &&
		(stq_valids_1[4] && stq_committed_1[4] ? !soc1.lsu._GEN_37481 : 1'b1) &&
		(stq_valids_1[5] && stq_committed_1[5] ? !soc1.lsu._GEN_37482 : 1'b1) &&
		(stq_valids_1[6] && stq_committed_1[6] ? !soc1.lsu._GEN_37483 : 1'b1) &&
		(stq_valids_1[7] && stq_committed_1[7] ? !soc1.lsu._GEN_37484 : 1'b1) &&
		(stq_valids_1[8] && stq_committed_1[8] ? !soc1.lsu._GEN_37485 : 1'b1) &&
		(stq_valids_1[9] && stq_committed_1[9] ? !soc1.lsu._GEN_37486 : 1'b1) &&
		(stq_valids_1[10] && stq_committed_1[10] ? !soc1.lsu._GEN_37487 : 1'b1) &&
		(stq_valids_1[11] && stq_committed_1[11] ? !soc1.lsu._GEN_37488 : 1'b1) &&
		(stq_valids_1[12] && stq_committed_1[12] ? !soc1.lsu._GEN_37489 : 1'b1) &&
		(stq_valids_1[13] && stq_committed_1[13] ? !soc1.lsu._GEN_37490 : 1'b1) &&
		(stq_valids_1[14] && stq_committed_1[14] ? !soc1.lsu._GEN_37491 : 1'b1) &&
		(stq_valids_1[15] && stq_committed_1[15] ? !soc1.lsu._GEN_37492 : 1'b1);
		
	wire exe_reg_0_sfence_not_speculative_1;
	assign exe_reg_0_sfence_not_speculative_1 = soc1.core.iregister_read.exe_reg_valids_0 && soc1.core.iregister_read.exe_reg_uops_0_mem_cmd == 5'h14 ? soc1.core.iregister_read.exe_reg_uops_0_br_mask == 12'h0 : 1'b1; 
	
	wire rrd_no_rocc_1;
	assign rrd_no_rocc_1 =
	(soc1.core.iregister_read.rrd_uops_0_REG_uopc != 7'h6c) && (soc1.core.iregister_read.rrd_uops_1_REG_uopc != 7'h6c) && (soc1.core.iregister_read.rrd_uops_2_REG_uopc != 7'h6c);
	
	wire dmem_req_amo_1;
	assign dmem_req_amo_1 = soc1.lsu.io_dmem_req_bits_0_valid && soc1.lsu.io_dmem_req_bits_0_bits_uop_is_amo? soc1.lsu.io_dmem_req_bits_0_bits_uop_br_mask == 12'h0 : 1'b1;
	
	wire fpu_req_uopc_1;
	assign fpu_req_uopc_1 = !soc1.core.fp_pipeline.fpiu_unit.fpu.io_req_valid || check_fpu_uopc(soc1.core.fp_pipeline.fpiu_unit.fpu.io_req_bits_uop_uopc);

	function automatic check_fpu_uopc(input [6:0] uopc);
	begin
	  case (uopc)
	    7'h48 : check_fpu_uopc = 1'b1; // uopFSGNJ_S
	    7'h49 : check_fpu_uopc = 1'b1; // uopFSGNJ_D
	    7'h4a : check_fpu_uopc = 1'b1; // uopFCVT_S_D
	    7'h4b : check_fpu_uopc = 1'b1; // uopFCVT_D_S
	    7'h54 : check_fpu_uopc = 1'b1; // uopFMINMAX_S
	    7'h55 : check_fpu_uopc = 1'b1; // uopFMINMAX_D
	    7'h57 : check_fpu_uopc = 1'b1; // uopFADD_S
	    7'h58 : check_fpu_uopc = 1'b1; // uopFSUB_S
	    7'h59 : check_fpu_uopc = 1'b1; // uopFMUL_S
	    7'h5a : check_fpu_uopc = 1'b1; // uopFADD_D
	    7'h5b : check_fpu_uopc = 1'b1; // uopFSUB_D
	    7'h5c : check_fpu_uopc = 1'b1; // uopFMUL_D
	    7'h5d : check_fpu_uopc = 1'b1; // uopFMADD_S
	    7'h5e : check_fpu_uopc = 1'b1; // uopFMSUB_S
	    7'h5f : check_fpu_uopc = 1'b1; // uopFNMADD_S
	    7'h60 : check_fpu_uopc = 1'b1; // uopFNMSUB_S
	    7'h61 : check_fpu_uopc = 1'b1; // uopFMADD_D
	    7'h62 : check_fpu_uopc = 1'b1; // uopFMSUB_D
	    7'h63 : check_fpu_uopc = 1'b1; // uopFNMADD_D
	    7'h64 : check_fpu_uopc = 1'b1; // uopFNMSUB_D
	    7'h52 : check_fpu_uopc = 1'b1; // uopFCLASS_S
	    7'h53 : check_fpu_uopc = 1'b1; // uopFCLASS_D
	    7'h46 : check_fpu_uopc = 1'b1; // uopFMV_X_S
	    7'h47 : check_fpu_uopc = 1'b1; // uopFMV_X_D
	    7'h4e : check_fpu_uopc = 1'b1; // uopFCVT_X_S
	    7'h4f : check_fpu_uopc = 1'b1; // uopFCVT_X_D
	    7'h50 : check_fpu_uopc = 1'b1; // uopCMPR_S
    	    7'h51 : check_fpu_uopc = 1'b1; // uopCMPR_D
    	    7'h2  : check_fpu_uopc = 1'b1; // uopSTA
	    default : check_fpu_uopc = 1'b0;
	  endcase
	end
	endfunction
	
	wire fdivsqrt_req_uopc_1;
	assign fdivsqrt_req_uopc_1 = !soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.io_req_valid || check_fdivsqrt_uopc(soc1.core.fp_pipeline.fpiu_unit.fdivsqrt.io_req_bits_uop_uopc);

	function automatic check_fdivsqrt_uopc(input [6:0] uopc);
	begin
	  case (uopc)
	    7'h65 : check_fdivsqrt_uopc = 1'b1; // uopFDIV_S
	    7'h66 : check_fdivsqrt_uopc = 1'b1; // uopFDIV_D
	    7'h67 : check_fdivsqrt_uopc = 1'b1; // uopFSQRT_S
	    7'h68 : check_fdivsqrt_uopc = 1'b1; // uopFSQRT_D
	    default : check_fdivsqrt_uopc = 1'b0;
	  endcase
	end
	endfunction
	
	wire fp_sdq_req_uopc_1;
	assign fp_sdq_req_uopc_1 = !soc1.core.fp_pipeline.fpiu_unit.fp_sdq.io_enq_valid || soc1.core.fp_pipeline.fpiu_unit.fp_sdq.io_enq_bits_uop_uopc == 7'h2;
	
	wire jmp_unit_ifpu_req_uopc_1;
	assign jmp_unit_ifpu_req_uopc_1 = !soc1.core.jmp_unit.ifpu.io_req_valid || check_jmp_unit_ifpu_uopc(soc1.core.jmp_unit.ifpu.io_req_bits_uop_uopc);

	function automatic check_jmp_unit_ifpu_uopc(input [6:0] uopc);
	begin
	  case (uopc)
	    7'h44 : check_jmp_unit_ifpu_uopc = 1'b1; // uopFMV_S_X
	    7'h45 : check_jmp_unit_ifpu_uopc = 1'b1; // uopFMV_D_X
	    7'h4c : check_jmp_unit_ifpu_uopc = 1'b1; // uopFCVT_S_X
	    7'h4d : check_jmp_unit_ifpu_uopc = 1'b1; // uopFCVT_D_X
	    default : check_jmp_unit_ifpu_uopc = 1'b0;
	  endcase
	end
	endfunction
	
	wire br_jal_jalr_consistent_uopc_1;
	assign br_jal_jalr_consistent_uopc_1 =
	(soc1.core.iregister_read.exe_reg_uops_1_is_br
	?
		soc1.core.iregister_read.exe_reg_uops_1_uopc == 7'h18 || soc1.core.iregister_read.exe_reg_uops_1_uopc == 7'h19 || soc1.core.iregister_read.exe_reg_uops_1_uopc == 7'h1a ||
		soc1.core.iregister_read.exe_reg_uops_1_uopc == 7'h1b || soc1.core.iregister_read.exe_reg_uops_1_uopc == 7'h1c || soc1.core.iregister_read.exe_reg_uops_1_uopc == 7'h1d
	: 1'b1) &&
	(soc1.core.iregister_read.exe_reg_uops_1_is_jal ? soc1.core.iregister_read.exe_reg_uops_1_uopc == 7'h25 : 1'b1) &&
	(soc1.core.iregister_read.exe_reg_uops_1_is_jalr ? soc1.core.iregister_read.exe_reg_uops_1_uopc == 7'h26 : 1'b1) &&
	(soc1.core.iregister_read.exe_reg_uops_2_is_br
	?
		soc1.core.iregister_read.exe_reg_uops_2_uopc == 7'h18 || soc1.core.iregister_read.exe_reg_uops_2_uopc == 7'h19 || soc1.core.iregister_read.exe_reg_uops_2_uopc == 7'h1a ||
		soc1.core.iregister_read.exe_reg_uops_2_uopc == 7'h1b || soc1.core.iregister_read.exe_reg_uops_2_uopc == 7'h1c || soc1.core.iregister_read.exe_reg_uops_2_uopc == 7'h1d
	: 1'b1) &&
	(soc1.core.iregister_read.exe_reg_uops_2_is_jal ? soc1.core.iregister_read.exe_reg_uops_2_uopc == 7'h25 : 1'b1) &&
	(soc1.core.iregister_read.exe_reg_uops_2_is_jalr ? soc1.core.iregister_read.exe_reg_uops_2_uopc == 7'h26 : 1'b1);

	//br_type and uopc consistent
	wire br_type_consistent_1;
	assign br_type_consistent_1 =
		(soc1.core.iregister_read.exe_reg_uops_1_ctrl_br_type == 4'h8 ? soc1.core.iregister_read.exe_reg_uops_1_uopc == 7'h26 : 1'b1) &&
    		(soc1.core.iregister_read.exe_reg_uops_2_ctrl_br_type == 4'h8 ? soc1.core.iregister_read.exe_reg_uops_2_uopc == 7'h26 : 1'b1);
    	    
    	wire sfence_at_head_1;
    	assign sfence_at_head_1 =
    		soc1.core.mem_units_0.maddrcalc.io_resp_bits_sfence_valid ? soc1.core.mem_units_0.maddrcalc.io_resp_bits_uop_rob_idx == soc1.core.rob.io_rob_head_idx : 1'b1;
	
	//wire ifpu_valids_consistent_1;
	//assign ifpu_valids_consistent_1 = soc1.core.jmp_unit.ifpu.ifpu.io_out_v ? soc1.core.jmp_unit.ifpu.r_valids_1 : 1'b1;
	
	//SoC2

  	//Create an array of the branch masks of the ROB
	wire [11:0] rob_branch_masks_2 [63:0];
	assign rob_branch_masks_2[0] = soc2.core.rob.rob_uop__0_br_mask;
	assign rob_branch_masks_2[1] = soc2.core.rob.rob_uop_1_0_br_mask;
	assign rob_branch_masks_2[2] = soc2.core.rob.rob_uop__1_br_mask;
	assign rob_branch_masks_2[3] = soc2.core.rob.rob_uop_1_1_br_mask;
	assign rob_branch_masks_2[4] = soc2.core.rob.rob_uop__2_br_mask;
	assign rob_branch_masks_2[5] = soc2.core.rob.rob_uop_1_2_br_mask;
	assign rob_branch_masks_2[6] = soc2.core.rob.rob_uop__3_br_mask;
	assign rob_branch_masks_2[7] = soc2.core.rob.rob_uop_1_3_br_mask;
	assign rob_branch_masks_2[8] = soc2.core.rob.rob_uop__4_br_mask;
	assign rob_branch_masks_2[9] = soc2.core.rob.rob_uop_1_4_br_mask;
	assign rob_branch_masks_2[10] = soc2.core.rob.rob_uop__5_br_mask;
	assign rob_branch_masks_2[11] = soc2.core.rob.rob_uop_1_5_br_mask;
	assign rob_branch_masks_2[12] = soc2.core.rob.rob_uop__6_br_mask;
	assign rob_branch_masks_2[13] = soc2.core.rob.rob_uop_1_6_br_mask;
	assign rob_branch_masks_2[14] = soc2.core.rob.rob_uop__7_br_mask;
	assign rob_branch_masks_2[15] = soc2.core.rob.rob_uop_1_7_br_mask;
	assign rob_branch_masks_2[16] = soc2.core.rob.rob_uop__8_br_mask;
	assign rob_branch_masks_2[17] = soc2.core.rob.rob_uop_1_8_br_mask;
	assign rob_branch_masks_2[18] = soc2.core.rob.rob_uop__9_br_mask;
	assign rob_branch_masks_2[19] = soc2.core.rob.rob_uop_1_9_br_mask;
	assign rob_branch_masks_2[20] = soc2.core.rob.rob_uop__10_br_mask;
	assign rob_branch_masks_2[21] = soc2.core.rob.rob_uop_1_10_br_mask;
	assign rob_branch_masks_2[22] = soc2.core.rob.rob_uop__11_br_mask;
	assign rob_branch_masks_2[23] = soc2.core.rob.rob_uop_1_11_br_mask;
	assign rob_branch_masks_2[24] = soc2.core.rob.rob_uop__12_br_mask;
	assign rob_branch_masks_2[25] = soc2.core.rob.rob_uop_1_12_br_mask;
	assign rob_branch_masks_2[26] = soc2.core.rob.rob_uop__13_br_mask;
	assign rob_branch_masks_2[27] = soc2.core.rob.rob_uop_1_13_br_mask;
	assign rob_branch_masks_2[28] = soc2.core.rob.rob_uop__14_br_mask;
	assign rob_branch_masks_2[29] = soc2.core.rob.rob_uop_1_14_br_mask;
	assign rob_branch_masks_2[30] = soc2.core.rob.rob_uop__15_br_mask;
	assign rob_branch_masks_2[31] = soc2.core.rob.rob_uop_1_15_br_mask;
	assign rob_branch_masks_2[32] = soc2.core.rob.rob_uop__16_br_mask;
	assign rob_branch_masks_2[33] = soc2.core.rob.rob_uop_1_16_br_mask;
	assign rob_branch_masks_2[34] = soc2.core.rob.rob_uop__17_br_mask;
	assign rob_branch_masks_2[35] = soc2.core.rob.rob_uop_1_17_br_mask;
	assign rob_branch_masks_2[36] = soc2.core.rob.rob_uop__18_br_mask;
	assign rob_branch_masks_2[37] = soc2.core.rob.rob_uop_1_18_br_mask;
	assign rob_branch_masks_2[38] = soc2.core.rob.rob_uop__19_br_mask;
	assign rob_branch_masks_2[39] = soc2.core.rob.rob_uop_1_19_br_mask;
	assign rob_branch_masks_2[40] = soc2.core.rob.rob_uop__20_br_mask;
	assign rob_branch_masks_2[41] = soc2.core.rob.rob_uop_1_20_br_mask;
	assign rob_branch_masks_2[42] = soc2.core.rob.rob_uop__21_br_mask;
	assign rob_branch_masks_2[43] = soc2.core.rob.rob_uop_1_21_br_mask;
	assign rob_branch_masks_2[44] = soc2.core.rob.rob_uop__22_br_mask;
	assign rob_branch_masks_2[45] = soc2.core.rob.rob_uop_1_22_br_mask;
	assign rob_branch_masks_2[46] = soc2.core.rob.rob_uop__23_br_mask;
	assign rob_branch_masks_2[47] = soc2.core.rob.rob_uop_1_23_br_mask;
	assign rob_branch_masks_2[48] = soc2.core.rob.rob_uop__24_br_mask;
	assign rob_branch_masks_2[49] = soc2.core.rob.rob_uop_1_24_br_mask;
	assign rob_branch_masks_2[50] = soc2.core.rob.rob_uop__25_br_mask;
	assign rob_branch_masks_2[51] = soc2.core.rob.rob_uop_1_25_br_mask;
	assign rob_branch_masks_2[52] = soc2.core.rob.rob_uop__26_br_mask;
	assign rob_branch_masks_2[53] = soc2.core.rob.rob_uop_1_26_br_mask;
	assign rob_branch_masks_2[54] = soc2.core.rob.rob_uop__27_br_mask;
	assign rob_branch_masks_2[55] = soc2.core.rob.rob_uop_1_27_br_mask;
	assign rob_branch_masks_2[56] = soc2.core.rob.rob_uop__28_br_mask;
	assign rob_branch_masks_2[57] = soc2.core.rob.rob_uop_1_28_br_mask;
	assign rob_branch_masks_2[58] = soc2.core.rob.rob_uop__29_br_mask;
	assign rob_branch_masks_2[59] = soc2.core.rob.rob_uop_1_29_br_mask;
	assign rob_branch_masks_2[60] = soc2.core.rob.rob_uop__30_br_mask;
	assign rob_branch_masks_2[61] = soc2.core.rob.rob_uop_1_30_br_mask;
	assign rob_branch_masks_2[62] = soc2.core.rob.rob_uop__31_br_mask;
	assign rob_branch_masks_2[63] = soc2.core.rob.rob_uop_1_31_br_mask;

	//Create an array of the valid bits of the ROB
	wire rob_valids_2 [63:0];
	assign rob_valids_2[0] = soc2.core.rob.rob_val__0;
	assign rob_valids_2[1] = soc2.core.rob.rob_val_1_0;
	assign rob_valids_2[2] = soc2.core.rob.rob_val__1;
	assign rob_valids_2[3] = soc2.core.rob.rob_val_1_1;
	assign rob_valids_2[4] = soc2.core.rob.rob_val__2;
	assign rob_valids_2[5] = soc2.core.rob.rob_val_1_2;
	assign rob_valids_2[6] = soc2.core.rob.rob_val__3;
	assign rob_valids_2[7] = soc2.core.rob.rob_val_1_3;
	assign rob_valids_2[8] = soc2.core.rob.rob_val__4;
	assign rob_valids_2[9] = soc2.core.rob.rob_val_1_4;
	assign rob_valids_2[10] = soc2.core.rob.rob_val__5;
	assign rob_valids_2[11] = soc2.core.rob.rob_val_1_5;
	assign rob_valids_2[12] = soc2.core.rob.rob_val__6;
	assign rob_valids_2[13] = soc2.core.rob.rob_val_1_6;
	assign rob_valids_2[14] = soc2.core.rob.rob_val__7;
	assign rob_valids_2[15] = soc2.core.rob.rob_val_1_7;
	assign rob_valids_2[16] = soc2.core.rob.rob_val__8;
	assign rob_valids_2[17] = soc2.core.rob.rob_val_1_8;
	assign rob_valids_2[18] = soc2.core.rob.rob_val__9;
	assign rob_valids_2[19] = soc2.core.rob.rob_val_1_9;
	assign rob_valids_2[20] = soc2.core.rob.rob_val__10;
	assign rob_valids_2[21] = soc2.core.rob.rob_val_1_10;
	assign rob_valids_2[22] = soc2.core.rob.rob_val__11;
	assign rob_valids_2[23] = soc2.core.rob.rob_val_1_11;
	assign rob_valids_2[24] = soc2.core.rob.rob_val__12;
	assign rob_valids_2[25] = soc2.core.rob.rob_val_1_12;
	assign rob_valids_2[26] = soc2.core.rob.rob_val__13;
	assign rob_valids_2[27] = soc2.core.rob.rob_val_1_13;
	assign rob_valids_2[28] = soc2.core.rob.rob_val__14;
	assign rob_valids_2[29] = soc2.core.rob.rob_val_1_14;
	assign rob_valids_2[30] = soc2.core.rob.rob_val__15;
	assign rob_valids_2[31] = soc2.core.rob.rob_val_1_15;
	assign rob_valids_2[32] = soc2.core.rob.rob_val__16;
	assign rob_valids_2[33] = soc2.core.rob.rob_val_1_16;
	assign rob_valids_2[34] = soc2.core.rob.rob_val__17;
	assign rob_valids_2[35] = soc2.core.rob.rob_val_1_17;
	assign rob_valids_2[36] = soc2.core.rob.rob_val__18;
	assign rob_valids_2[37] = soc2.core.rob.rob_val_1_18;
	assign rob_valids_2[38] = soc2.core.rob.rob_val__19;
	assign rob_valids_2[39] = soc2.core.rob.rob_val_1_19;
	assign rob_valids_2[40] = soc2.core.rob.rob_val__20;
	assign rob_valids_2[41] = soc2.core.rob.rob_val_1_20;
	assign rob_valids_2[42] = soc2.core.rob.rob_val__21;
	assign rob_valids_2[43] = soc2.core.rob.rob_val_1_21;
	assign rob_valids_2[44] = soc2.core.rob.rob_val__22;
	assign rob_valids_2[45] = soc2.core.rob.rob_val_1_22;
	assign rob_valids_2[46] = soc2.core.rob.rob_val__23;
	assign rob_valids_2[47] = soc2.core.rob.rob_val_1_23;
	assign rob_valids_2[48] = soc2.core.rob.rob_val__24;
	assign rob_valids_2[49] = soc2.core.rob.rob_val_1_24;
	assign rob_valids_2[50] = soc2.core.rob.rob_val__25;
	assign rob_valids_2[51] = soc2.core.rob.rob_val_1_25;
	assign rob_valids_2[52] = soc2.core.rob.rob_val__26;
	assign rob_valids_2[53] = soc2.core.rob.rob_val_1_26;
	assign rob_valids_2[54] = soc2.core.rob.rob_val__27;
	assign rob_valids_2[55] = soc2.core.rob.rob_val_1_27;
	assign rob_valids_2[56] = soc2.core.rob.rob_val__28;
	assign rob_valids_2[57] = soc2.core.rob.rob_val_1_28;
	assign rob_valids_2[58] = soc2.core.rob.rob_val__29;
	assign rob_valids_2[59] = soc2.core.rob.rob_val_1_29;
	assign rob_valids_2[60] = soc2.core.rob.rob_val__30;
	assign rob_valids_2[61] = soc2.core.rob.rob_val_1_30;
	assign rob_valids_2[62] = soc2.core.rob.rob_val__31;
	assign rob_valids_2[63] = soc2.core.rob.rob_val_1_31;

	//array that stores a copy of the rob_idx of the ldq
	wire [5:0] ldq_rob_idx_2 [15:0];
	assign ldq_rob_idx_2[0] = soc2.lsu.ldq_0_bits_uop_rob_idx;
	assign ldq_rob_idx_2[1] = soc2.lsu.ldq_1_bits_uop_rob_idx;
	assign ldq_rob_idx_2[2] = soc2.lsu.ldq_2_bits_uop_rob_idx;
	assign ldq_rob_idx_2[3] = soc2.lsu.ldq_3_bits_uop_rob_idx;
	assign ldq_rob_idx_2[4] = soc2.lsu.ldq_4_bits_uop_rob_idx;
	assign ldq_rob_idx_2[5] = soc2.lsu.ldq_5_bits_uop_rob_idx;
	assign ldq_rob_idx_2[6] = soc2.lsu.ldq_6_bits_uop_rob_idx;
	assign ldq_rob_idx_2[7] = soc2.lsu.ldq_7_bits_uop_rob_idx;
	assign ldq_rob_idx_2[8] = soc2.lsu.ldq_8_bits_uop_rob_idx;
	assign ldq_rob_idx_2[9] = soc2.lsu.ldq_9_bits_uop_rob_idx;
	assign ldq_rob_idx_2[10] = soc2.lsu.ldq_10_bits_uop_rob_idx;
	assign ldq_rob_idx_2[11] = soc2.lsu.ldq_11_bits_uop_rob_idx;
	assign ldq_rob_idx_2[12] = soc2.lsu.ldq_12_bits_uop_rob_idx;
	assign ldq_rob_idx_2[13] = soc2.lsu.ldq_13_bits_uop_rob_idx;
	assign ldq_rob_idx_2[14] = soc2.lsu.ldq_14_bits_uop_rob_idx;
	assign ldq_rob_idx_2[15] = soc2.lsu.ldq_15_bits_uop_rob_idx;

	wire rob_uses_stq_2 [63:0];
	assign rob_uses_stq_2[0] = soc2.core.rob.rob_uop__0_uses_stq;
	assign rob_uses_stq_2[1] = soc2.core.rob.rob_uop_1_0_uses_stq;
	assign rob_uses_stq_2[2] = soc2.core.rob.rob_uop__1_uses_stq;
	assign rob_uses_stq_2[3] = soc2.core.rob.rob_uop_1_1_uses_stq;
	assign rob_uses_stq_2[4] = soc2.core.rob.rob_uop__2_uses_stq;
	assign rob_uses_stq_2[5] = soc2.core.rob.rob_uop_1_2_uses_stq;
	assign rob_uses_stq_2[6] = soc2.core.rob.rob_uop__3_uses_stq;
	assign rob_uses_stq_2[7] = soc2.core.rob.rob_uop_1_3_uses_stq;
	assign rob_uses_stq_2[8] = soc2.core.rob.rob_uop__4_uses_stq;
	assign rob_uses_stq_2[9] = soc2.core.rob.rob_uop_1_4_uses_stq;
	assign rob_uses_stq_2[10] = soc2.core.rob.rob_uop__5_uses_stq;
	assign rob_uses_stq_2[11] = soc2.core.rob.rob_uop_1_5_uses_stq;
	assign rob_uses_stq_2[12] = soc2.core.rob.rob_uop__6_uses_stq;
	assign rob_uses_stq_2[13] = soc2.core.rob.rob_uop_1_6_uses_stq;
	assign rob_uses_stq_2[14] = soc2.core.rob.rob_uop__7_uses_stq;
	assign rob_uses_stq_2[15] = soc2.core.rob.rob_uop_1_7_uses_stq;
	assign rob_uses_stq_2[16] = soc2.core.rob.rob_uop__8_uses_stq;
	assign rob_uses_stq_2[17] = soc2.core.rob.rob_uop_1_8_uses_stq;
	assign rob_uses_stq_2[18] = soc2.core.rob.rob_uop__9_uses_stq;
	assign rob_uses_stq_2[19] = soc2.core.rob.rob_uop_1_9_uses_stq;
	assign rob_uses_stq_2[20] = soc2.core.rob.rob_uop__10_uses_stq;
	assign rob_uses_stq_2[21] = soc2.core.rob.rob_uop_1_10_uses_stq;
	assign rob_uses_stq_2[22] = soc2.core.rob.rob_uop__11_uses_stq;
	assign rob_uses_stq_2[23] = soc2.core.rob.rob_uop_1_11_uses_stq;
	assign rob_uses_stq_2[24] = soc2.core.rob.rob_uop__12_uses_stq;
	assign rob_uses_stq_2[25] = soc2.core.rob.rob_uop_1_12_uses_stq;
	assign rob_uses_stq_2[26] = soc2.core.rob.rob_uop__13_uses_stq;
	assign rob_uses_stq_2[27] = soc2.core.rob.rob_uop_1_13_uses_stq;
	assign rob_uses_stq_2[28] = soc2.core.rob.rob_uop__14_uses_stq;
	assign rob_uses_stq_2[29] = soc2.core.rob.rob_uop_1_14_uses_stq;
	assign rob_uses_stq_2[30] = soc2.core.rob.rob_uop__15_uses_stq;
	assign rob_uses_stq_2[31] = soc2.core.rob.rob_uop_1_15_uses_stq;
	assign rob_uses_stq_2[32] = soc2.core.rob.rob_uop__16_uses_stq;
	assign rob_uses_stq_2[33] = soc2.core.rob.rob_uop_1_16_uses_stq;
	assign rob_uses_stq_2[34] = soc2.core.rob.rob_uop__17_uses_stq;
	assign rob_uses_stq_2[35] = soc2.core.rob.rob_uop_1_17_uses_stq;
	assign rob_uses_stq_2[36] = soc2.core.rob.rob_uop__18_uses_stq;
	assign rob_uses_stq_2[37] = soc2.core.rob.rob_uop_1_18_uses_stq;
	assign rob_uses_stq_2[38] = soc2.core.rob.rob_uop__19_uses_stq;
	assign rob_uses_stq_2[39] = soc2.core.rob.rob_uop_1_19_uses_stq;
	assign rob_uses_stq_2[40] = soc2.core.rob.rob_uop__20_uses_stq;
	assign rob_uses_stq_2[41] = soc2.core.rob.rob_uop_1_20_uses_stq;
	assign rob_uses_stq_2[42] = soc2.core.rob.rob_uop__21_uses_stq;
	assign rob_uses_stq_2[43] = soc2.core.rob.rob_uop_1_21_uses_stq;
	assign rob_uses_stq_2[44] = soc2.core.rob.rob_uop__22_uses_stq;
	assign rob_uses_stq_2[45] = soc2.core.rob.rob_uop_1_22_uses_stq;
	assign rob_uses_stq_2[46] = soc2.core.rob.rob_uop__23_uses_stq;
	assign rob_uses_stq_2[47] = soc2.core.rob.rob_uop_1_23_uses_stq;
	assign rob_uses_stq_2[48] = soc2.core.rob.rob_uop__24_uses_stq;
	assign rob_uses_stq_2[49] = soc2.core.rob.rob_uop_1_24_uses_stq;
	assign rob_uses_stq_2[50] = soc2.core.rob.rob_uop__25_uses_stq;
	assign rob_uses_stq_2[51] = soc2.core.rob.rob_uop_1_25_uses_stq;
	assign rob_uses_stq_2[52] = soc2.core.rob.rob_uop__26_uses_stq;
	assign rob_uses_stq_2[53] = soc2.core.rob.rob_uop_1_26_uses_stq;
	assign rob_uses_stq_2[54] = soc2.core.rob.rob_uop__27_uses_stq;
	assign rob_uses_stq_2[55] = soc2.core.rob.rob_uop_1_27_uses_stq;
	assign rob_uses_stq_2[56] = soc2.core.rob.rob_uop__28_uses_stq;
	assign rob_uses_stq_2[57] = soc2.core.rob.rob_uop_1_28_uses_stq;
	assign rob_uses_stq_2[58] = soc2.core.rob.rob_uop__29_uses_stq;
	assign rob_uses_stq_2[59] = soc2.core.rob.rob_uop_1_29_uses_stq;
	assign rob_uses_stq_2[60] = soc2.core.rob.rob_uop__30_uses_stq;
	assign rob_uses_stq_2[61] = soc2.core.rob.rob_uop_1_30_uses_stq;
	assign rob_uses_stq_2[62] = soc2.core.rob.rob_uop__31_uses_stq;
	assign rob_uses_stq_2[63] = soc2.core.rob.rob_uop_1_31_uses_stq;

	wire rob_uses_ldq_2 [63:0];
	assign rob_uses_ldq_2[0] = soc2.core.rob.rob_uop__0_uses_ldq;
	assign rob_uses_ldq_2[1] = soc2.core.rob.rob_uop_1_0_uses_ldq;
	assign rob_uses_ldq_2[2] = soc2.core.rob.rob_uop__1_uses_ldq;
	assign rob_uses_ldq_2[3] = soc2.core.rob.rob_uop_1_1_uses_ldq;
	assign rob_uses_ldq_2[4] = soc2.core.rob.rob_uop__2_uses_ldq;
	assign rob_uses_ldq_2[5] = soc2.core.rob.rob_uop_1_2_uses_ldq;
	assign rob_uses_ldq_2[6] = soc2.core.rob.rob_uop__3_uses_ldq;
	assign rob_uses_ldq_2[7] = soc2.core.rob.rob_uop_1_3_uses_ldq;
	assign rob_uses_ldq_2[8] = soc2.core.rob.rob_uop__4_uses_ldq;
	assign rob_uses_ldq_2[9] = soc2.core.rob.rob_uop_1_4_uses_ldq;
	assign rob_uses_ldq_2[10] = soc2.core.rob.rob_uop__5_uses_ldq;
	assign rob_uses_ldq_2[11] = soc2.core.rob.rob_uop_1_5_uses_ldq;
	assign rob_uses_ldq_2[12] = soc2.core.rob.rob_uop__6_uses_ldq;
	assign rob_uses_ldq_2[13] = soc2.core.rob.rob_uop_1_6_uses_ldq;
	assign rob_uses_ldq_2[14] = soc2.core.rob.rob_uop__7_uses_ldq;
	assign rob_uses_ldq_2[15] = soc2.core.rob.rob_uop_1_7_uses_ldq;
	assign rob_uses_ldq_2[16] = soc2.core.rob.rob_uop__8_uses_ldq;
	assign rob_uses_ldq_2[17] = soc2.core.rob.rob_uop_1_8_uses_ldq;
	assign rob_uses_ldq_2[18] = soc2.core.rob.rob_uop__9_uses_ldq;
	assign rob_uses_ldq_2[19] = soc2.core.rob.rob_uop_1_9_uses_ldq;
	assign rob_uses_ldq_2[20] = soc2.core.rob.rob_uop__10_uses_ldq;
	assign rob_uses_ldq_2[21] = soc2.core.rob.rob_uop_1_10_uses_ldq;
	assign rob_uses_ldq_2[22] = soc2.core.rob.rob_uop__11_uses_ldq;
	assign rob_uses_ldq_2[23] = soc2.core.rob.rob_uop_1_11_uses_ldq;
	assign rob_uses_ldq_2[24] = soc2.core.rob.rob_uop__12_uses_ldq;
	assign rob_uses_ldq_2[25] = soc2.core.rob.rob_uop_1_12_uses_ldq;
	assign rob_uses_ldq_2[26] = soc2.core.rob.rob_uop__13_uses_ldq;
	assign rob_uses_ldq_2[27] = soc2.core.rob.rob_uop_1_13_uses_ldq;
	assign rob_uses_ldq_2[28] = soc2.core.rob.rob_uop__14_uses_ldq;
	assign rob_uses_ldq_2[29] = soc2.core.rob.rob_uop_1_14_uses_ldq;
	assign rob_uses_ldq_2[30] = soc2.core.rob.rob_uop__15_uses_ldq;
	assign rob_uses_ldq_2[31] = soc2.core.rob.rob_uop_1_15_uses_ldq;
	assign rob_uses_ldq_2[32] = soc2.core.rob.rob_uop__16_uses_ldq;
	assign rob_uses_ldq_2[33] = soc2.core.rob.rob_uop_1_16_uses_ldq;
	assign rob_uses_ldq_2[34] = soc2.core.rob.rob_uop__17_uses_ldq;
	assign rob_uses_ldq_2[35] = soc2.core.rob.rob_uop_1_17_uses_ldq;
	assign rob_uses_ldq_2[36] = soc2.core.rob.rob_uop__18_uses_ldq;
	assign rob_uses_ldq_2[37] = soc2.core.rob.rob_uop_1_18_uses_ldq;
	assign rob_uses_ldq_2[38] = soc2.core.rob.rob_uop__19_uses_ldq;
	assign rob_uses_ldq_2[39] = soc2.core.rob.rob_uop_1_19_uses_ldq;
	assign rob_uses_ldq_2[40] = soc2.core.rob.rob_uop__20_uses_ldq;
	assign rob_uses_ldq_2[41] = soc2.core.rob.rob_uop_1_20_uses_ldq;
	assign rob_uses_ldq_2[42] = soc2.core.rob.rob_uop__21_uses_ldq;
	assign rob_uses_ldq_2[43] = soc2.core.rob.rob_uop_1_21_uses_ldq;
	assign rob_uses_ldq_2[44] = soc2.core.rob.rob_uop__22_uses_ldq;
	assign rob_uses_ldq_2[45] = soc2.core.rob.rob_uop_1_22_uses_ldq;
	assign rob_uses_ldq_2[46] = soc2.core.rob.rob_uop__23_uses_ldq;
	assign rob_uses_ldq_2[47] = soc2.core.rob.rob_uop_1_23_uses_ldq;
	assign rob_uses_ldq_2[48] = soc2.core.rob.rob_uop__24_uses_ldq;
	assign rob_uses_ldq_2[49] = soc2.core.rob.rob_uop_1_24_uses_ldq;
	assign rob_uses_ldq_2[50] = soc2.core.rob.rob_uop__25_uses_ldq;
	assign rob_uses_ldq_2[51] = soc2.core.rob.rob_uop_1_25_uses_ldq;
	assign rob_uses_ldq_2[52] = soc2.core.rob.rob_uop__26_uses_ldq;
	assign rob_uses_ldq_2[53] = soc2.core.rob.rob_uop_1_26_uses_ldq;
	assign rob_uses_ldq_2[54] = soc2.core.rob.rob_uop__27_uses_ldq;
	assign rob_uses_ldq_2[55] = soc2.core.rob.rob_uop_1_27_uses_ldq;
	assign rob_uses_ldq_2[56] = soc2.core.rob.rob_uop__28_uses_ldq;
	assign rob_uses_ldq_2[57] = soc2.core.rob.rob_uop_1_28_uses_ldq;
	assign rob_uses_ldq_2[58] = soc2.core.rob.rob_uop__29_uses_ldq;
	assign rob_uses_ldq_2[59] = soc2.core.rob.rob_uop_1_29_uses_ldq;
	assign rob_uses_ldq_2[60] = soc2.core.rob.rob_uop__30_uses_ldq;
	assign rob_uses_ldq_2[61] = soc2.core.rob.rob_uop_1_30_uses_ldq;
	assign rob_uses_ldq_2[62] = soc2.core.rob.rob_uop__31_uses_ldq;
	assign rob_uses_ldq_2[63] = soc2.core.rob.rob_uop_1_31_uses_ldq;
	
	//Create an array of the exception bits of the ROB
	wire rob_exception_2 [63:0];
	assign rob_exception_2[0] = soc2.core.rob.rob_exception__0;
	assign rob_exception_2[1] = soc2.core.rob.rob_exception_1_0;
	assign rob_exception_2[2] = soc2.core.rob.rob_exception__1;
	assign rob_exception_2[3] = soc2.core.rob.rob_exception_1_1;
	assign rob_exception_2[4] = soc2.core.rob.rob_exception__2;
	assign rob_exception_2[5] = soc2.core.rob.rob_exception_1_2;
	assign rob_exception_2[6] = soc2.core.rob.rob_exception__3;
	assign rob_exception_2[7] = soc2.core.rob.rob_exception_1_3;
	assign rob_exception_2[8] = soc2.core.rob.rob_exception__4;
	assign rob_exception_2[9] = soc2.core.rob.rob_exception_1_4;
	assign rob_exception_2[10] = soc2.core.rob.rob_exception__5;
	assign rob_exception_2[11] = soc2.core.rob.rob_exception_1_5;
	assign rob_exception_2[12] = soc2.core.rob.rob_exception__6;
	assign rob_exception_2[13] = soc2.core.rob.rob_exception_1_6;
	assign rob_exception_2[14] = soc2.core.rob.rob_exception__7;
	assign rob_exception_2[15] = soc2.core.rob.rob_exception_1_7;
	assign rob_exception_2[16] = soc2.core.rob.rob_exception__8;
	assign rob_exception_2[17] = soc2.core.rob.rob_exception_1_8;
	assign rob_exception_2[18] = soc2.core.rob.rob_exception__9;
	assign rob_exception_2[19] = soc2.core.rob.rob_exception_1_9;
	assign rob_exception_2[20] = soc2.core.rob.rob_exception__10;
	assign rob_exception_2[21] = soc2.core.rob.rob_exception_1_10;
	assign rob_exception_2[22] = soc2.core.rob.rob_exception__11;
	assign rob_exception_2[23] = soc2.core.rob.rob_exception_1_11;
	assign rob_exception_2[24] = soc2.core.rob.rob_exception__12;
	assign rob_exception_2[25] = soc2.core.rob.rob_exception_1_12;
	assign rob_exception_2[26] = soc2.core.rob.rob_exception__13;
	assign rob_exception_2[27] = soc2.core.rob.rob_exception_1_13;
	assign rob_exception_2[28] = soc2.core.rob.rob_exception__14;
	assign rob_exception_2[29] = soc2.core.rob.rob_exception_1_14;
	assign rob_exception_2[30] = soc2.core.rob.rob_exception__15;
	assign rob_exception_2[31] = soc2.core.rob.rob_exception_1_15;
	assign rob_exception_2[32] = soc2.core.rob.rob_exception__16;
	assign rob_exception_2[33] = soc2.core.rob.rob_exception_1_16;
	assign rob_exception_2[34] = soc2.core.rob.rob_exception__17;
	assign rob_exception_2[35] = soc2.core.rob.rob_exception_1_17;
	assign rob_exception_2[36] = soc2.core.rob.rob_exception__18;
	assign rob_exception_2[37] = soc2.core.rob.rob_exception_1_18;
	assign rob_exception_2[38] = soc2.core.rob.rob_exception__19;
	assign rob_exception_2[39] = soc2.core.rob.rob_exception_1_19;
	assign rob_exception_2[40] = soc2.core.rob.rob_exception__20;
	assign rob_exception_2[41] = soc2.core.rob.rob_exception_1_20;
	assign rob_exception_2[42] = soc2.core.rob.rob_exception__21;
	assign rob_exception_2[43] = soc2.core.rob.rob_exception_1_21;
	assign rob_exception_2[44] = soc2.core.rob.rob_exception__22;
	assign rob_exception_2[45] = soc2.core.rob.rob_exception_1_22;
	assign rob_exception_2[46] = soc2.core.rob.rob_exception__23;
	assign rob_exception_2[47] = soc2.core.rob.rob_exception_1_23;
	assign rob_exception_2[48] = soc2.core.rob.rob_exception__24;
	assign rob_exception_2[49] = soc2.core.rob.rob_exception_1_24;
	assign rob_exception_2[50] = soc2.core.rob.rob_exception__25;
	assign rob_exception_2[51] = soc2.core.rob.rob_exception_1_25;
	assign rob_exception_2[52] = soc2.core.rob.rob_exception__26;
	assign rob_exception_2[53] = soc2.core.rob.rob_exception_1_26;
	assign rob_exception_2[54] = soc2.core.rob.rob_exception__27;
	assign rob_exception_2[55] = soc2.core.rob.rob_exception_1_27;
	assign rob_exception_2[56] = soc2.core.rob.rob_exception__28;
	assign rob_exception_2[57] = soc2.core.rob.rob_exception_1_28;
	assign rob_exception_2[58] = soc2.core.rob.rob_exception__29;
	assign rob_exception_2[59] = soc2.core.rob.rob_exception_1_29;
	assign rob_exception_2[60] = soc2.core.rob.rob_exception__30;
	assign rob_exception_2[61] = soc2.core.rob.rob_exception_1_30;
	assign rob_exception_2[62] = soc2.core.rob.rob_exception__31;
	assign rob_exception_2[63] = soc2.core.rob.rob_exception_1_31;

	//array that stores a copy of the rob_idx of the stq
	wire [5:0] stq_rob_idx_2 [15:0];
	assign stq_rob_idx_2[0] = soc2.lsu.stq_0_bits_uop_rob_idx;
	assign stq_rob_idx_2[1] = soc2.lsu.stq_1_bits_uop_rob_idx;
	assign stq_rob_idx_2[2] = soc2.lsu.stq_2_bits_uop_rob_idx;
	assign stq_rob_idx_2[3] = soc2.lsu.stq_3_bits_uop_rob_idx;
	assign stq_rob_idx_2[4] = soc2.lsu.stq_4_bits_uop_rob_idx;
	assign stq_rob_idx_2[5] = soc2.lsu.stq_5_bits_uop_rob_idx;
	assign stq_rob_idx_2[6] = soc2.lsu.stq_6_bits_uop_rob_idx;
	assign stq_rob_idx_2[7] = soc2.lsu.stq_7_bits_uop_rob_idx;
	assign stq_rob_idx_2[8] = soc2.lsu.stq_8_bits_uop_rob_idx;
	assign stq_rob_idx_2[9] = soc2.lsu.stq_9_bits_uop_rob_idx;
	assign stq_rob_idx_2[10] = soc2.lsu.stq_10_bits_uop_rob_idx;
	assign stq_rob_idx_2[11] = soc2.lsu.stq_11_bits_uop_rob_idx;
	assign stq_rob_idx_2[12] = soc2.lsu.stq_12_bits_uop_rob_idx;
	assign stq_rob_idx_2[13] = soc2.lsu.stq_13_bits_uop_rob_idx;
	assign stq_rob_idx_2[14] = soc2.lsu.stq_14_bits_uop_rob_idx;
	assign stq_rob_idx_2[15] = soc2.lsu.stq_15_bits_uop_rob_idx;

	//array that stores a copy of the committed bits of the stq
	wire stq_committed_2 [15:0];
	assign stq_committed_2[0] = soc2.lsu.stq_0_bits_committed;
	assign stq_committed_2[1] = soc2.lsu.stq_1_bits_committed;
	assign stq_committed_2[2] = soc2.lsu.stq_2_bits_committed;
	assign stq_committed_2[3] = soc2.lsu.stq_3_bits_committed;
	assign stq_committed_2[4] = soc2.lsu.stq_4_bits_committed;
	assign stq_committed_2[5] = soc2.lsu.stq_5_bits_committed;
	assign stq_committed_2[6] = soc2.lsu.stq_6_bits_committed;
	assign stq_committed_2[7] = soc2.lsu.stq_7_bits_committed;
	assign stq_committed_2[8] = soc2.lsu.stq_8_bits_committed;
	assign stq_committed_2[9] = soc2.lsu.stq_9_bits_committed;
	assign stq_committed_2[10] = soc2.lsu.stq_10_bits_committed;
	assign stq_committed_2[11] = soc2.lsu.stq_11_bits_committed;
	assign stq_committed_2[12] = soc2.lsu.stq_12_bits_committed;
	assign stq_committed_2[13] = soc2.lsu.stq_13_bits_committed;
	assign stq_committed_2[14] = soc2.lsu.stq_14_bits_committed;
	assign stq_committed_2[15] = soc2.lsu.stq_15_bits_committed;

	//function that returns true if the given ID in ROB is above or equal ldq_head and below ldq_tail
	function automatic isInBoundsROB_2;
	  //6-bit ID of the ROB entry
	  input [5:0] id;
	  begin
	    if(rob_valids_2[id] == 1'b1)
	    begin
	      //distinguish between positions of head and tail
	      if (soc2.core.rob.io_rob_head_idx < soc2.core.rob.io_rob_tail_idx)
	      begin
	  isInBoundsROB_2 = (id >= soc2.core.rob.io_rob_head_idx && id < soc2.core.rob.io_rob_tail_idx) || soc2.core.rob.full;
	      end
	      else if (soc2.core.rob.io_rob_head_idx > soc2.core.rob.io_rob_tail_idx)
	      begin
	  isInBoundsROB_2 = (id >= soc2.core.rob.io_rob_head_idx || id < soc2.core.rob.io_rob_tail_idx) || soc2.core.rob.full;
	      end
	      else // soc2.core.rob.io_rob_head_idx == soc2.core.rob.io_rob_tail_idx
	      begin
	  isInBoundsROB_2 = !soc2.core.rob.io_empty;
	      end
	    end
	    else
	    begin
	      isInBoundsROB_2 = 1'b0;
	    end
	  end
	endfunction

  wire consistent_branch_masks_2;
	assign consistent_branch_masks_2 =
	(
	//is the uop at head valid and is the ROB not empty
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 0) % 64)
	?
	  (
	  //if true, the branch mask at head must be 0 because the first valid instruction after head must be non-speculative
	  rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 0) % 64] == 12'b0
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 1) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 0) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 0) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 1) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 0) % 64]
	  :
	    (
	    //if head is invalid, the branch mask at head + 1 must be 0 because the first valid instruction after head must be non-speculative
	    rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] == 12'b0
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 2) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 2) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 1) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 0) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 0) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 2) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 0) % 64]
	    :
	      //if head is invalid, the branch mask at head + 2 must be 0 because the first valid instruction after head must be non-speculative
	      rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] == 12'b0
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 3) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 3) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 2) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 3) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 1) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 0) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 3) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 0) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 4) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 4) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 3) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 4) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 2) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 4) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 1) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 5) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 5) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 4) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 5) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 3) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 5) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 2) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 6) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 6) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 5) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 6) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 4) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 6) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 3) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 7) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 7) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 6) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 7) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 5) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 7) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 4) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 8) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 8) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 7) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 8) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 6) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 8) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 5) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 9) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 9) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 8) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 9) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 7) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 9) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 6) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 10) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 10) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 9) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 10) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 8) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 10) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 7) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 11) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 11) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 10) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 11) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 9) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 11) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 8) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 12) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 12) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 11) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 12) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 10) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 12) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 9) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 13) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 13) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 12) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 13) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 11) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 13) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 10) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 14) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 14) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 13) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 14) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 12) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 14) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 11) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 15) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 15) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 14) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 15) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 13) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 15) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 12) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 16) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 16) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 15) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 16) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 14) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 16) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 13) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 17) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 17) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 16) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 17) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 15) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 17) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 14) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 18) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 18) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 17) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 18) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 16) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 18) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 15) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 19) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 19) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 18) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 19) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 17) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 19) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 16) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 20) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 20) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 19) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 20) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 18) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 20) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 17) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 21) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 21) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 20) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 21) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 19) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 21) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 18) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 22) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 22) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 21) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 22) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 20) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 22) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 19) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 23) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 23) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 22) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 23) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 21) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 23) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 20) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 24) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 24) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 23) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 24) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 22) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 24) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 21) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 25) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 25) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 24) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 25) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 23) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 25) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 22) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 26) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 26) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 25) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 26) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 24) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 26) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 23) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 27) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 27) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 26) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 27) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 25) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 27) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 24) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 28) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 28) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 27) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 28) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 26) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 28) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 25) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 29) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 29) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 28) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 29) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 27) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 29) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 26) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 30) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 30) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 29) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 30) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 28) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 30) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 27) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 31) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 31) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 30) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 31) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 29) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 31) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 28) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 32) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 32) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 31) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 32) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 30) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 32) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 29) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 33) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 33) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 32) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 33) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 31) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 33) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 30) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 34) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 34) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 33) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 34) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 32) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 34) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 31) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 35) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 35) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 34) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 35) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 33) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 35) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 32) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 36) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 36) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 35) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 36) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 34) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 36) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 33) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 37) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 37) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 36) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 37) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 35) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 37) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 34) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 38) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 38) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 37) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 38) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 36) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 38) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 35) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 39) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 39) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 38) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 39) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 37) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 39) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 36) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 40) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 40) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 39) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 40) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 38) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 40) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 37) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 41) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 41) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 40) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 41) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 39) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 41) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 38) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 42) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 42) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 41) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 42) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 40) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 42) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 39) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 43) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 43) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 42) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 43) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 41) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 43) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 40) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 44) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 44) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 43) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 44) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 42) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 44) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 41) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 45) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 45) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 44) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 45) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 43) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 45) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 42) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 46) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 46) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 45) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 46) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 44) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 46) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 43) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 47) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 47) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 46) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 47) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 45) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 47) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 44) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 48) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 48) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 47) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 48) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 46) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 48) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 45) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 49) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 49) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 48) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 49) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 47) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 49) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 46) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 50) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 50) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 49) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 50) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 48) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 50) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 47) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 51) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 51) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 50) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 51) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 49) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 51) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 48) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 52) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 52) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 51) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 52) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 50) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 52) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 49) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 53) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 53) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 52) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 53) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 51) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 53) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 50) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 54) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 54) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 53) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 54) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 52) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 54) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 51) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 55) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 55) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 54) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 55) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 53) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 55) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 52) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 56) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 56) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 55) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 56) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 54) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 56) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 53) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 57) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 57) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 56) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 57) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 55) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 57) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 54) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 58) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 58) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 57) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 58) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 56) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 58) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 55) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 59) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 59) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 58) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 59) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 57) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 59) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 56) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 60) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 60) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 59) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 60) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 58) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 60) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 57) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 61) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 61) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 60) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 61) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 59) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 61) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 58) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 62) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 61) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 62) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 61) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 62) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 60) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 62) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 59) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	) &&
	(
	//is the uop at head + X in between head and tail and is it valid?
	isInBoundsROB_2((soc2.core.rob.io_rob_head_idx + 63) % 64)
	?
	  (
	  //check if the prior uop X-1 is a valid one
	  rob_valids_2[(soc2.core.rob.io_rob_head_idx + 62) % 64] == 1'b1
	  ?
	    // do a bitwise AND on the branch masks of uop X and X-1
	    // this has to be equal to the branch mask of X-1
	    (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 62) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 63) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 62) % 64]
	  :
	    (
	    //in case X-1 is a bubble/invalid instruction
	    //go another step back to X-2 and check its validity
	    rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64] == 1'b1
	    ?
	      //compare branch masks of X and X-2 then
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 61) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 63) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 61) % 64]
	    :
	      //else compare with X-3 (there SHOULD not be any empty rows, so at least X-3 has to be valid)
	      (rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] & rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 63) % 64]) == rob_branch_masks_2[(soc2.core.rob.io_rob_head_idx + 60) % 64]
	    )
	  )
	:
	  //else branch mask can be arbitrary
	  1'b1
	);

	wire consistent_valid_flags_2;
	assign consistent_valid_flags_2 =
	(
	soc2.core.rob.io_empty == 1'b1
	?
		//if empty, no entry can be valid
		(soc2.core.rob.rob_val__0 | soc2.core.rob.rob_val_1_0 | soc2.core.rob.rob_val__1 | soc2.core.rob.rob_val_1_1 | soc2.core.rob.rob_val__2 | soc2.core.rob.rob_val_1_2 |
		soc2.core.rob.rob_val__3 | soc2.core.rob.rob_val_1_3 | soc2.core.rob.rob_val__4 | soc2.core.rob.rob_val_1_4 | soc2.core.rob.rob_val__5 | soc2.core.rob.rob_val_1_5 |
		soc2.core.rob.rob_val__6 | soc2.core.rob.rob_val_1_6 | soc2.core.rob.rob_val__7 | soc2.core.rob.rob_val_1_7 | soc2.core.rob.rob_val__8 | soc2.core.rob.rob_val_1_8 |
		soc2.core.rob.rob_val__9 | soc2.core.rob.rob_val_1_9 | soc2.core.rob.rob_val__10 | soc2.core.rob.rob_val_1_10 | soc2.core.rob.rob_val__11 | soc2.core.rob.rob_val_1_11 |
		soc2.core.rob.rob_val__12 | soc2.core.rob.rob_val_1_12 | soc2.core.rob.rob_val__13 | soc2.core.rob.rob_val_1_13 | soc2.core.rob.rob_val__14 | soc2.core.rob.rob_val_1_14 |
		soc2.core.rob.rob_val__15 | soc2.core.rob.rob_val_1_15 | soc2.core.rob.rob_val__16 | soc2.core.rob.rob_val_1_16 | soc2.core.rob.rob_val__17 | soc2.core.rob.rob_val_1_17 |
		soc2.core.rob.rob_val__18 | soc2.core.rob.rob_val_1_18 | soc2.core.rob.rob_val__19 | soc2.core.rob.rob_val_1_19 | soc2.core.rob.rob_val__20 | soc2.core.rob.rob_val_1_20 |
		soc2.core.rob.rob_val__21 | soc2.core.rob.rob_val_1_21 | soc2.core.rob.rob_val__22 | soc2.core.rob.rob_val_1_22 | soc2.core.rob.rob_val__23 | soc2.core.rob.rob_val_1_23 |
		soc2.core.rob.rob_val__24 | soc2.core.rob.rob_val_1_24 | soc2.core.rob.rob_val__25 | soc2.core.rob.rob_val_1_25 | soc2.core.rob.rob_val__26 | soc2.core.rob.rob_val_1_26 |
		soc2.core.rob.rob_val__27 | soc2.core.rob.rob_val_1_27 | soc2.core.rob.rob_val__28 | soc2.core.rob.rob_val_1_28 | soc2.core.rob.rob_val__29 | soc2.core.rob.rob_val_1_29 |
		soc2.core.rob.rob_val__30 | soc2.core.rob.rob_val_1_30 | soc2.core.rob.rob_val__31 | soc2.core.rob.rob_val_1_31) == 1'b0
	:
		//if not empty
		//check for branch misprediction
		soc2.core.b2_mispredict
		?
			//only entries that are older than the mispredicted branch and the mispredicted branch itself can be valid
			//distinction for different head_lsbs
			(soc2.core.rob.rob_head_lsb == 1'b0)
			?
				//if not empty, at least one entry at head is valid
				//check for every entry if it is older than b2_uop_rob_idx + 1
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 0) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 0) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 0) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 1) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 0) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 1) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 2) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 2) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 4) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 4) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 6) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 6) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 8) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 8) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 10) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 10) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 12) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 12) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 14) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 14) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 16) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 16) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 18) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 18) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 20) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 20) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 22) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 22) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 24) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 24) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 26) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 26) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 28) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 28) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 30) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 30) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 32) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 32) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 34) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 34) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 36) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 36) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 38) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 38) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 40) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 40) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 42) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 42) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 44) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 44) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 46) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 46) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 48) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 48) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 50) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 50) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 52) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 52) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 54) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 54) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 56) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 56) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 58) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 58) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 60) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 60) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 62) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 62) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 62) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 63) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 62) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 63) % 64])
				)
			:
				//else if rob_head_lsb==1'b1
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 0) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 0) % 64) == soc2.core.b2_uop_rob_idx
				? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 0) % 64]
				: !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 0) % 64]
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 1) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 1) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 3) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 3) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 5) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 5) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 7) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 7) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 9) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 9) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 11) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 11) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 13) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 13) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 15) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 15) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 17) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 17) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 19) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 19) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 21) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 21) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 23) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 23) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 25) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 25) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 27) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 27) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 29) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 29) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 31) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 31) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 33) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 33) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 35) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 35) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 37) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 37) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 39) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 39) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 41) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 41) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 43) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 43) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 45) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 45) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 47) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 47) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 49) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 49) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 51) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 51) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 53) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 53) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 55) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 55) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 57) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 57) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 59) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 59) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 61) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 61) % 64) == soc2.core.b2_uop_rob_idx
				? (rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 62) % 64])
				: (!rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 62) % 64])
				) &&
				(ROBisOlder((soc2.core.rob.io_rob_head_idx + 63) % 64, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) || ((soc2.core.rob.io_rob_head_idx + 63) % 64) == soc2.core.b2_uop_rob_idx
				? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 63) % 64]
				: !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 63) % 64]
				)
		:
			soc2.core.rob.full == 1'b1
			?
				//if full, at least one entry per row has to be valid
				(soc2.core.rob.rob_val__0 || soc2.core.rob.rob_val_1_0) && (soc2.core.rob.rob_val__1 || soc2.core.rob.rob_val_1_1) && (soc2.core.rob.rob_val__2 || soc2.core.rob.rob_val_1_2) &&
				(soc2.core.rob.rob_val__3 || soc2.core.rob.rob_val_1_3) && (soc2.core.rob.rob_val__4 || soc2.core.rob.rob_val_1_4) && (soc2.core.rob.rob_val__5 || soc2.core.rob.rob_val_1_5) &&
				(soc2.core.rob.rob_val__6 || soc2.core.rob.rob_val_1_6) && (soc2.core.rob.rob_val__7 || soc2.core.rob.rob_val_1_7) && (soc2.core.rob.rob_val__8 || soc2.core.rob.rob_val_1_8) &&
				(soc2.core.rob.rob_val__9 || soc2.core.rob.rob_val_1_9) && (soc2.core.rob.rob_val__10 || soc2.core.rob.rob_val_1_10) && (soc2.core.rob.rob_val__11 || soc2.core.rob.rob_val_1_11) &&
				(soc2.core.rob.rob_val__12 || soc2.core.rob.rob_val_1_12) && (soc2.core.rob.rob_val__13 || soc2.core.rob.rob_val_1_13) && (soc2.core.rob.rob_val__14 || soc2.core.rob.rob_val_1_14) &&
				(soc2.core.rob.rob_val__15 || soc2.core.rob.rob_val_1_15) && (soc2.core.rob.rob_val__16 || soc2.core.rob.rob_val_1_16) && (soc2.core.rob.rob_val__17 || soc2.core.rob.rob_val_1_17) &&
				(soc2.core.rob.rob_val__18 || soc2.core.rob.rob_val_1_18) && (soc2.core.rob.rob_val__19 || soc2.core.rob.rob_val_1_19) && (soc2.core.rob.rob_val__20 || soc2.core.rob.rob_val_1_20) &&
				(soc2.core.rob.rob_val__21 || soc2.core.rob.rob_val_1_21) && (soc2.core.rob.rob_val__22 || soc2.core.rob.rob_val_1_22) && (soc2.core.rob.rob_val__23 || soc2.core.rob.rob_val_1_23) &&
				(soc2.core.rob.rob_val__24 || soc2.core.rob.rob_val_1_24) && (soc2.core.rob.rob_val__25 || soc2.core.rob.rob_val_1_25) && (soc2.core.rob.rob_val__26 || soc2.core.rob.rob_val_1_26) &&
				(soc2.core.rob.rob_val__27 || soc2.core.rob.rob_val_1_27) && (soc2.core.rob.rob_val__28 || soc2.core.rob.rob_val_1_28) && (soc2.core.rob.rob_val__29 || soc2.core.rob.rob_val_1_29) &&
				(soc2.core.rob.rob_val__30 || soc2.core.rob.rob_val_1_30) && (soc2.core.rob.rob_val__31 || soc2.core.rob.rob_val_1_31)
			:
				//if not empty, full, rollback or branch mispredict
				//in every row, that is older than tail there has to be at least one valid entry
				//distinction for different head_lsbs
				(
				(soc2.core.rob.rob_head_lsb == 1'b0)
				?
					//if neither full or empty, at least one entry at head is valid
					(rob_valids_2[(soc2.core.rob.io_rob_head_idx + 0) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 1) % 64]) &&
					//for every row that is before tail, there is at least one valid entry
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 2) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 4) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 6) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 8) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 10) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 12) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 14) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 16) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 18) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 20) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 22) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 24) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 26) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 28) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 30) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 32) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 34) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 36) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 38) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 40) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 42) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 44) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 46) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 48) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 50) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 52) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 54) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 56) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 58) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 60) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 62) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 62) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 63) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 62) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 63) % 64]) &&
					//make sure that tail points an invalid entry
					(soc2.core.rob.rob_state == 2'h2 ? 1'b1 : rob_valids_2[soc2.core.rob.io_rob_tail_idx] == 1'b0)
				:
					//if soc2.core.rob.rob_head_lsb == 1'b1
					//if neither full or empty, head must be valid, since head_lsb is 1
					(rob_valids_2[(soc2.core.rob.io_rob_head_idx + 0) % 64]) &&
					//for every row that is before tail, there is at least one valid entry
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 1) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 1) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 2) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 3) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 3) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 4) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 5) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 5) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 6) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 7) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 7) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 8) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 9) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 9) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 10) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 11) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 11) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 12) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 13) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 13) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 14) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 15) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 15) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 16) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 17) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 17) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 18) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 19) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 19) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 20) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 21) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 21) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 22) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 23) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 23) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 24) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 25) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 25) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 26) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 27) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 27) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 28) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 29) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 29) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 30) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 31) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 31) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 32) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 33) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 33) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 34) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 35) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 35) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 36) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 37) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 37) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 38) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 39) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 39) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 40) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 41) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 41) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 42) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 43) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 43) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 44) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 45) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 45) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 46) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 47) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 47) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 48) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 49) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 49) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 50) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 51) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 51) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 52) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 53) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 53) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 54) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 55) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 55) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 56) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 57) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 57) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 58) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 59) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 59) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 60) % 64]) &&
					((ROBisOlder((soc2.core.rob.io_rob_head_idx + 61) % 64, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx)) ? rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64] || rob_valids_2[(soc2.core.rob.io_rob_head_idx + 62) % 64] : !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 61) % 64] && !rob_valids_2[(soc2.core.rob.io_rob_head_idx + 62) % 64]) &&
					//head+63 is in fact the entry before head+0, which must be invalid, since ROB is not full
					(rob_valids_2[(soc2.core.rob.io_rob_head_idx + 63) % 64] == 1'b0) &&
					//make sure that tail points an invalid entry
					(soc2.core.rob.rob_state == 2'h2 ? 1'b1 : rob_valids_2[soc2.core.rob.io_rob_tail_idx] == 1'b0)
				)
	);



	//if tail is rolled back because of a mispredict, make sure it is rolled back to an older value than tail
	wire consistent_tail_rollback_2;
	assign consistent_tail_rollback_2 =
	  (soc2.core.b2_mispredict == 1'b1 ? ROBisOlder(soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx) || soc2.core.rob.full: 1'b1)
	;

	//ensure that no speculative instruction commits
	wire no_speculative_commit_2;
	assign no_speculative_commit_2 =
	  (soc2.core.rob.will_commit_0 ? (rob_branch_masks_2[{soc2.core.rob.rob_head, 1'b0}] == 12'b0) && rob_branch_masks_2[soc2.core.rob.io_commit_uops_0_rob_idx] == 12'b0 : 1'b1) &&
	  (soc2.core.rob.will_commit_1 ? (rob_branch_masks_2[{soc2.core.rob.rob_head, 1'b1}] == 12'b0) && rob_branch_masks_2[soc2.core.rob.io_commit_uops_0_rob_idx] == 12'b0 : 1'b1)
	;

	//function that returns true if the given ID in store queue is above or equal stq_head and below stq_tail
	function automatic isInBoundsSTQ_2;
	//4-bit ID of the store queue entry
	input [3:0] id;
	begin
	//distinguish between positions of head and tail
	if (soc2.lsu.stq_head < soc2.lsu.stq_tail)
	begin
	  isInBoundsSTQ_2 =  id >= soc2.lsu.stq_head && id < soc2.lsu.stq_tail;
	end
	else if (soc2.lsu.stq_head > soc2.lsu.stq_tail)
	begin
	  isInBoundsSTQ_2 = id >= soc2.lsu.stq_head || id < soc2.lsu.stq_tail;
	end
	else // soc2.lsu.stq_head == soc2.lsu.stq_tail
	begin
	  isInBoundsSTQ_2 = 1'b1; // stq is full or empty, handled separately
	end
	end
	endfunction

	//stores that are not inside FIFO bounds have to be invalid to avoid unreachable dependencies
	wire stq_check_invalidated_entries_2;
	assign stq_check_invalidated_entries_2 =
	//check if misprediction happened last cycle
	  (soc2.core.b2_mispredict
	    ?
	    (isInBoundsSTQ_2(4'h0) && ROBisOlder(soc2.lsu.stq_0_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_0_valid : !soc2.lsu.stq_0_valid || soc2.lsu.stq_0_bits_committed) &&
	    (isInBoundsSTQ_2(4'h1) && ROBisOlder(soc2.lsu.stq_1_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_1_valid : !soc2.lsu.stq_1_valid || soc2.lsu.stq_1_bits_committed) &&
	    (isInBoundsSTQ_2(4'h2) && ROBisOlder(soc2.lsu.stq_2_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_2_valid : !soc2.lsu.stq_2_valid || soc2.lsu.stq_2_bits_committed) &&
	    (isInBoundsSTQ_2(4'h3) && ROBisOlder(soc2.lsu.stq_3_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_3_valid : !soc2.lsu.stq_3_valid || soc2.lsu.stq_3_bits_committed) &&
	    (isInBoundsSTQ_2(4'h4) && ROBisOlder(soc2.lsu.stq_4_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_4_valid : !soc2.lsu.stq_4_valid || soc2.lsu.stq_4_bits_committed) &&
	    (isInBoundsSTQ_2(4'h5) && ROBisOlder(soc2.lsu.stq_5_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_5_valid : !soc2.lsu.stq_5_valid || soc2.lsu.stq_5_bits_committed) &&
	    (isInBoundsSTQ_2(4'h6) && ROBisOlder(soc2.lsu.stq_6_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_6_valid : !soc2.lsu.stq_6_valid || soc2.lsu.stq_6_bits_committed) &&
	    (isInBoundsSTQ_2(4'h7) && ROBisOlder(soc2.lsu.stq_7_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_7_valid : !soc2.lsu.stq_7_valid || soc2.lsu.stq_7_bits_committed) &&
	    (isInBoundsSTQ_2(4'h8) && ROBisOlder(soc2.lsu.stq_8_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_8_valid : !soc2.lsu.stq_8_valid || soc2.lsu.stq_8_bits_committed) &&
	    (isInBoundsSTQ_2(4'h9) && ROBisOlder(soc2.lsu.stq_9_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_9_valid : !soc2.lsu.stq_9_valid || soc2.lsu.stq_9_bits_committed) &&
	    (isInBoundsSTQ_2(4'ha) && ROBisOlder(soc2.lsu.stq_10_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_10_valid : !soc2.lsu.stq_10_valid || soc2.lsu.stq_10_bits_committed) &&
	    (isInBoundsSTQ_2(4'hb) && ROBisOlder(soc2.lsu.stq_11_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_11_valid : !soc2.lsu.stq_11_valid || soc2.lsu.stq_11_bits_committed) &&
	    (isInBoundsSTQ_2(4'hc) && ROBisOlder(soc2.lsu.stq_12_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_12_valid : !soc2.lsu.stq_12_valid || soc2.lsu.stq_12_bits_committed) &&
	    (isInBoundsSTQ_2(4'hd) && ROBisOlder(soc2.lsu.stq_13_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_13_valid : !soc2.lsu.stq_13_valid || soc2.lsu.stq_13_bits_committed) &&
	    (isInBoundsSTQ_2(4'he) && ROBisOlder(soc2.lsu.stq_14_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_14_valid : !soc2.lsu.stq_14_valid || soc2.lsu.stq_14_bits_committed) &&
	    (isInBoundsSTQ_2(4'hf) && ROBisOlder(soc2.lsu.stq_15_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.stq_15_valid : !soc2.lsu.stq_15_valid || soc2.lsu.stq_15_bits_committed)
	    :
				//check if stq is empty, full or none of both
				((soc2.lsu.stq_head == soc2.lsu.stq_tail)
				?
					(soc2.lsu.stq_0_valid | soc2.lsu.stq_1_valid | soc2.lsu.stq_2_valid | soc2.lsu.stq_3_valid | soc2.lsu.stq_4_valid | soc2.lsu.stq_5_valid |	soc2.lsu.stq_6_valid | soc2.lsu.stq_7_valid | soc2.lsu.stq_8_valid | soc2.lsu.stq_12_valid | soc2.lsu.stq_13_valid | soc2.lsu.stq_14_valid | soc2.lsu.stq_15_valid)
					 == 1'b1
					 ?
				 		//if one is valid, stq has to be full
						(soc2.lsu.stq_0_valid & soc2.lsu.stq_1_valid & soc2.lsu.stq_2_valid &
						soc2.lsu.stq_3_valid & soc2.lsu.stq_4_valid & soc2.lsu.stq_5_valid &
						soc2.lsu.stq_6_valid & soc2.lsu.stq_7_valid & soc2.lsu.stq_8_valid &
						soc2.lsu.stq_9_valid & soc2.lsu.stq_10_valid & soc2.lsu.stq_11_valid &
						soc2.lsu.stq_12_valid & soc2.lsu.stq_13_valid & soc2.lsu.stq_14_valid &
						soc2.lsu.stq_15_valid) == 1'b1
					 :
						//if equal stq is empty
						(soc2.lsu.stq_0_valid | soc2.lsu.stq_1_valid | soc2.lsu.stq_2_valid |
						soc2.lsu.stq_3_valid | soc2.lsu.stq_4_valid | soc2.lsu.stq_5_valid |
						soc2.lsu.stq_6_valid | soc2.lsu.stq_7_valid | soc2.lsu.stq_8_valid |
						soc2.lsu.stq_9_valid | soc2.lsu.stq_10_valid | soc2.lsu.stq_11_valid |
						soc2.lsu.stq_12_valid | soc2.lsu.stq_13_valid | soc2.lsu.stq_14_valid |
						soc2.lsu.stq_15_valid) == 1'b0
				:
					//if not empty and not full, only valid bits with ID greater equal head or less than tail are set
					(isInBoundsSTQ_2(4'h0) ? soc2.lsu.stq_0_valid : !soc2.lsu.stq_0_valid) &&
					(isInBoundsSTQ_2(4'h1) ? soc2.lsu.stq_1_valid : !soc2.lsu.stq_1_valid) &&
					(isInBoundsSTQ_2(4'h2) ? soc2.lsu.stq_2_valid : !soc2.lsu.stq_2_valid) &&
					(isInBoundsSTQ_2(4'h3) ? soc2.lsu.stq_3_valid : !soc2.lsu.stq_3_valid) &&
					(isInBoundsSTQ_2(4'h4) ? soc2.lsu.stq_4_valid : !soc2.lsu.stq_4_valid) &&
					(isInBoundsSTQ_2(4'h5) ? soc2.lsu.stq_5_valid : !soc2.lsu.stq_5_valid) &&
					(isInBoundsSTQ_2(4'h6) ? soc2.lsu.stq_6_valid : !soc2.lsu.stq_6_valid) &&
					(isInBoundsSTQ_2(4'h7) ? soc2.lsu.stq_7_valid : !soc2.lsu.stq_7_valid) &&
					(isInBoundsSTQ_2(4'h8) ? soc2.lsu.stq_8_valid : !soc2.lsu.stq_8_valid) &&
					(isInBoundsSTQ_2(4'h9) ? soc2.lsu.stq_9_valid : !soc2.lsu.stq_9_valid) &&
					(isInBoundsSTQ_2(4'ha) ? soc2.lsu.stq_10_valid : !soc2.lsu.stq_10_valid) &&
					(isInBoundsSTQ_2(4'hb) ? soc2.lsu.stq_11_valid : !soc2.lsu.stq_11_valid) &&
					(isInBoundsSTQ_2(4'hc) ? soc2.lsu.stq_12_valid : !soc2.lsu.stq_12_valid) &&
					(isInBoundsSTQ_2(4'hd) ? soc2.lsu.stq_13_valid : !soc2.lsu.stq_13_valid) &&
					(isInBoundsSTQ_2(4'he) ? soc2.lsu.stq_14_valid : !soc2.lsu.stq_14_valid) &&
					(isInBoundsSTQ_2(4'hf) ? soc2.lsu.stq_15_valid : !soc2.lsu.stq_15_valid)
	  			)
	);

	//function that returns true if the given ID in load queue is above or equal ldq_head and below ldq_tail
	function automatic isInBoundsLDQ_2;
	  //4-bit ID of the load queue entry
	  input [3:0] id;
	  begin
	    //distinguish between positions of head and tail
	    if (soc2.lsu.ldq_head < soc2.lsu.ldq_tail)
	    begin
	      isInBoundsLDQ_2 =  id >= soc2.lsu.ldq_head && id < soc2.lsu.ldq_tail;
	    end
	    else if (soc2.lsu.ldq_head > soc2.lsu.ldq_tail)
	    begin
	      isInBoundsLDQ_2 = id >= soc2.lsu.ldq_head || id < soc2.lsu.ldq_tail;
	    end
	    else // soc2.lsu.ldq_head == soc2.lsu.ldq_tail
	    begin
	      isInBoundsLDQ_2 = 1'b1; // ldq is full or empty, handled separately
	    end
	  end
	endfunction

	//loads that are not inside FIFO bounds have to be invalid to avoid unreachable dependencies
	wire ldq_check_invalidated_entries_2;
	assign ldq_check_invalidated_entries_2 =
	//check if misprediction happened last cycle
		soc2.core.b2_mispredict
		?
			(isInBoundsLDQ_2(4'h0) && ROBisOlder(soc2.lsu.ldq_0_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_0_valid : !soc2.lsu.ldq_0_valid) &&
			(isInBoundsLDQ_2(4'h1) && ROBisOlder(soc2.lsu.ldq_1_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_1_valid : !soc2.lsu.ldq_1_valid) &&
			(isInBoundsLDQ_2(4'h2) && ROBisOlder(soc2.lsu.ldq_2_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_2_valid : !soc2.lsu.ldq_2_valid) &&
			(isInBoundsLDQ_2(4'h3) && ROBisOlder(soc2.lsu.ldq_3_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_3_valid : !soc2.lsu.ldq_3_valid) &&
			(isInBoundsLDQ_2(4'h4) && ROBisOlder(soc2.lsu.ldq_4_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_4_valid : !soc2.lsu.ldq_4_valid) &&
			(isInBoundsLDQ_2(4'h5) && ROBisOlder(soc2.lsu.ldq_5_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_5_valid : !soc2.lsu.ldq_5_valid) &&
			(isInBoundsLDQ_2(4'h6) && ROBisOlder(soc2.lsu.ldq_6_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_6_valid : !soc2.lsu.ldq_6_valid) &&
			(isInBoundsLDQ_2(4'h7) && ROBisOlder(soc2.lsu.ldq_7_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_7_valid : !soc2.lsu.ldq_7_valid) &&
			(isInBoundsLDQ_2(4'h8) && ROBisOlder(soc2.lsu.ldq_8_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_8_valid : !soc2.lsu.ldq_8_valid) &&
			(isInBoundsLDQ_2(4'h9) && ROBisOlder(soc2.lsu.ldq_9_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_9_valid : !soc2.lsu.ldq_9_valid) &&
			(isInBoundsLDQ_2(4'ha) && ROBisOlder(soc2.lsu.ldq_10_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_10_valid : !soc2.lsu.ldq_10_valid) &&
			(isInBoundsLDQ_2(4'hb) && ROBisOlder(soc2.lsu.ldq_11_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_11_valid : !soc2.lsu.ldq_11_valid) &&
			(isInBoundsLDQ_2(4'hc) && ROBisOlder(soc2.lsu.ldq_12_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_12_valid : !soc2.lsu.ldq_12_valid) &&
			(isInBoundsLDQ_2(4'hd) && ROBisOlder(soc2.lsu.ldq_13_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_13_valid : !soc2.lsu.ldq_13_valid) &&
			(isInBoundsLDQ_2(4'he) && ROBisOlder(soc2.lsu.ldq_14_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_14_valid : !soc2.lsu.ldq_14_valid) &&
			(isInBoundsLDQ_2(4'hf) && ROBisOlder(soc2.lsu.ldq_15_bits_uop_rob_idx, soc2.core.b2_uop_rob_idx, soc2.core.rob.io_rob_head_idx) ? soc2.lsu.ldq_15_valid : !soc2.lsu.ldq_15_valid)
		:
			//if equal ldq is empty
			(soc2.lsu.ldq_head == soc2.lsu.ldq_tail
			?
		 		(soc2.lsu.ldq_0_valid | soc2.lsu.ldq_1_valid | soc2.lsu.ldq_2_valid | soc2.lsu.ldq_3_valid | soc2.lsu.ldq_4_valid | soc2.lsu.ldq_5_valid |	soc2.lsu.ldq_6_valid | soc2.lsu.ldq_7_valid | soc2.lsu.ldq_8_valid | soc2.lsu.ldq_12_valid | soc2.lsu.ldq_13_valid | soc2.lsu.ldq_14_valid | soc2.lsu.ldq_15_valid)
				 == 1'b1
				?
					//if one is valid, ldq has to be full
					(soc2.lsu.ldq_0_valid & soc2.lsu.ldq_1_valid & soc2.lsu.ldq_2_valid &
					soc2.lsu.ldq_3_valid & soc2.lsu.ldq_4_valid & soc2.lsu.ldq_5_valid &
					soc2.lsu.ldq_6_valid & soc2.lsu.ldq_7_valid & soc2.lsu.ldq_8_valid &
					soc2.lsu.ldq_9_valid & soc2.lsu.ldq_10_valid & soc2.lsu.ldq_11_valid &
					soc2.lsu.ldq_12_valid & soc2.lsu.ldq_13_valid & soc2.lsu.ldq_14_valid &
					soc2.lsu.ldq_15_valid) == 1'b1
				:
					//if empty all valid bits are zero
					(soc2.lsu.ldq_0_valid | soc2.lsu.ldq_1_valid | soc2.lsu.ldq_2_valid |
					soc2.lsu.ldq_3_valid | soc2.lsu.ldq_4_valid | soc2.lsu.ldq_5_valid |
					soc2.lsu.ldq_6_valid | soc2.lsu.ldq_7_valid | soc2.lsu.ldq_8_valid |
					soc2.lsu.ldq_9_valid | soc2.lsu.ldq_10_valid | soc2.lsu.ldq_11_valid |
					soc2.lsu.ldq_12_valid | soc2.lsu.ldq_13_valid | soc2.lsu.ldq_14_valid |
					soc2.lsu.ldq_15_valid) == 1'b0
			:
				//if not empty and not full, only valid bits with ID greater equal head or less than tail are set
				(isInBoundsLDQ_2(4'h0) ? soc2.lsu.ldq_0_valid : !soc2.lsu.ldq_0_valid) &&
				(isInBoundsLDQ_2(4'h1) ? soc2.lsu.ldq_1_valid : !soc2.lsu.ldq_1_valid) &&
				(isInBoundsLDQ_2(4'h2) ? soc2.lsu.ldq_2_valid : !soc2.lsu.ldq_2_valid) &&
				(isInBoundsLDQ_2(4'h3) ? soc2.lsu.ldq_3_valid : !soc2.lsu.ldq_3_valid) &&
				(isInBoundsLDQ_2(4'h4) ? soc2.lsu.ldq_4_valid : !soc2.lsu.ldq_4_valid) &&
				(isInBoundsLDQ_2(4'h5) ? soc2.lsu.ldq_5_valid : !soc2.lsu.ldq_5_valid) &&
				(isInBoundsLDQ_2(4'h6) ? soc2.lsu.ldq_6_valid : !soc2.lsu.ldq_6_valid) &&
				(isInBoundsLDQ_2(4'h7) ? soc2.lsu.ldq_7_valid : !soc2.lsu.ldq_7_valid) &&
				(isInBoundsLDQ_2(4'h8) ? soc2.lsu.ldq_8_valid : !soc2.lsu.ldq_8_valid) &&
				(isInBoundsLDQ_2(4'h9) ? soc2.lsu.ldq_9_valid : !soc2.lsu.ldq_9_valid) &&
				(isInBoundsLDQ_2(4'ha) ? soc2.lsu.ldq_10_valid : !soc2.lsu.ldq_10_valid) &&
				(isInBoundsLDQ_2(4'hb) ? soc2.lsu.ldq_11_valid : !soc2.lsu.ldq_11_valid) &&
				(isInBoundsLDQ_2(4'hc) ? soc2.lsu.ldq_12_valid : !soc2.lsu.ldq_12_valid) &&
				(isInBoundsLDQ_2(4'hd) ? soc2.lsu.ldq_13_valid : !soc2.lsu.ldq_13_valid) &&
				(isInBoundsLDQ_2(4'he) ? soc2.lsu.ldq_14_valid : !soc2.lsu.ldq_14_valid) &&
				(isInBoundsLDQ_2(4'hf) ? soc2.lsu.ldq_15_valid : !soc2.lsu.ldq_15_valid)
			)
	;

	wire consistent_buffer_br_masks_2;
	assign consistent_buffer_br_masks_2 =
	  (soc2.core.csr_exe_unit.alu.r_valids_0 ? rob_valids_2[soc2.core.csr_exe_unit.alu.r_uops_0_rob_idx] && soc2.core.csr_exe_unit.alu.r_uops_0_br_mask == rob_branch_masks_2[soc2.core.csr_exe_unit.alu.r_uops_0_rob_idx] : 1'b1) &&
	  ((soc2.core.csr_exe_unit.div.div.state == 3'h3) ||(soc2.core.csr_exe_unit.div.div.state == 3'h7) ? rob_valids_2[soc2.core.csr_exe_unit.div.r_uop_rob_idx] && soc2.core.csr_exe_unit.div.r_uop_br_mask == rob_branch_masks_2[soc2.core.csr_exe_unit.div.r_uop_rob_idx] : 1'b1) &&
	  (soc2.core.iregister_read.exe_reg_valids_0 /*&& !(soc2.core.iregister_read.exe_reg_uops_0_uses_stq && stq_committed_2[soc2.core.iregister_read.exe_reg_uops_0_stq_idx]) */? rob_valids_2[soc2.core.iregister_read.exe_reg_uops_0_rob_idx] && soc2.core.iregister_read.exe_reg_uops_0_br_mask == rob_branch_masks_2[soc2.core.iregister_read.exe_reg_uops_0_rob_idx] : 1'b1) &&
	  (soc2.core.iregister_read.exe_reg_valids_1 /*&& !(soc2.core.iregister_read.exe_reg_uops_1_uses_stq && stq_committed_2[soc2.core.iregister_read.exe_reg_uops_1_stq_idx]) */? rob_valids_2[soc2.core.iregister_read.exe_reg_uops_1_rob_idx] && soc2.core.iregister_read.exe_reg_uops_1_br_mask == rob_branch_masks_2[soc2.core.iregister_read.exe_reg_uops_1_rob_idx] : 1'b1) &&
	  (soc2.core.iregister_read.exe_reg_valids_2 /*&& !(soc2.core.iregister_read.exe_reg_uops_2_uses_stq && stq_committed_2[soc2.core.iregister_read.exe_reg_uops_2_stq_idx]) */? rob_valids_2[soc2.core.iregister_read.exe_reg_uops_2_rob_idx] && soc2.core.iregister_read.exe_reg_uops_2_br_mask == rob_branch_masks_2[soc2.core.iregister_read.exe_reg_uops_2_rob_idx] : 1'b1) &&
	  (soc2.core.iregister_read.rrd_valids_0_REG /*&& !(soc2.core.iregister_read.rrd_uops_0_REG_uses_stq && stq_committed_2[soc2.core.iregister_read.rrd_uops_0_REG_stq_idx]) */? rob_valids_2[soc2.core.iregister_read.rrd_uops_0_REG_rob_idx] && soc2.core.iregister_read.rrd_uops_0_REG_br_mask == rob_branch_masks_2[soc2.core.iregister_read.rrd_uops_0_REG_rob_idx] : 1'b1) &&
	  (soc2.core.iregister_read.rrd_valids_1_REG /*&& !(soc2.core.iregister_read.rrd_uops_1_REG_uses_stq && stq_committed_2[soc2.core.iregister_read.rrd_uops_1_REG_stq_idx]) */? rob_valids_2[soc2.core.iregister_read.rrd_uops_1_REG_rob_idx] && soc2.core.iregister_read.rrd_uops_1_REG_br_mask == rob_branch_masks_2[soc2.core.iregister_read.rrd_uops_1_REG_rob_idx] : 1'b1) &&
	  (soc2.core.iregister_read.rrd_valids_2_REG /*&& !(soc2.core.iregister_read.rrd_uops_2_REG_uses_stq && stq_committed_2[soc2.core.iregister_read.rrd_uops_2_REG_stq_idx]) */? rob_valids_2[soc2.core.iregister_read.rrd_uops_2_REG_rob_idx] && soc2.core.iregister_read.rrd_uops_2_REG_br_mask == rob_branch_masks_2[soc2.core.iregister_read.rrd_uops_2_REG_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.queue.valids_0 ? rob_valids_2[soc2.core.jmp_unit.queue.uops_0_rob_idx] && soc2.core.jmp_unit.queue.uops_0_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.queue.uops_0_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.queue.valids_1 ? rob_valids_2[soc2.core.jmp_unit.queue.uops_1_rob_idx] && soc2.core.jmp_unit.queue.uops_1_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.queue.uops_1_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.queue.valids_2 ? rob_valids_2[soc2.core.jmp_unit.queue.uops_2_rob_idx] && soc2.core.jmp_unit.queue.uops_2_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.queue.uops_2_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.queue.valids_3 ? rob_valids_2[soc2.core.jmp_unit.queue.uops_3_rob_idx] && soc2.core.jmp_unit.queue.uops_3_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.queue.uops_3_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.queue.valids_4 ? rob_valids_2[soc2.core.jmp_unit.queue.uops_4_rob_idx] && soc2.core.jmp_unit.queue.uops_4_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.queue.uops_4_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.alu.r_valids_0 ? rob_valids_2[soc2.core.jmp_unit.alu.r_uops_0_rob_idx] && soc2.core.jmp_unit.alu.r_uops_0_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.alu.r_uops_0_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.alu.r_valids_1 ? rob_valids_2[soc2.core.jmp_unit.alu.r_uops_1_rob_idx] && soc2.core.jmp_unit.alu.r_uops_1_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.alu.r_uops_1_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.alu.r_valids_2 ? rob_valids_2[soc2.core.jmp_unit.alu.r_uops_2_rob_idx] && soc2.core.jmp_unit.alu.r_uops_2_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.alu.r_uops_2_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.ifpu.r_valids_0 ? rob_valids_2[soc2.core.jmp_unit.ifpu.r_uops_0_rob_idx] && soc2.core.jmp_unit.ifpu.r_uops_0_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.ifpu.r_uops_0_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.ifpu.r_valids_1 ? rob_valids_2[soc2.core.jmp_unit.ifpu.r_uops_1_rob_idx] && soc2.core.jmp_unit.ifpu.r_uops_1_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.ifpu.r_uops_1_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.imul.r_valids_0 ? rob_valids_2[soc2.core.jmp_unit.imul.r_uops_0_rob_idx] && soc2.core.jmp_unit.imul.r_uops_0_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.imul.r_uops_0_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.imul.r_valids_1 ? rob_valids_2[soc2.core.jmp_unit.imul.r_uops_1_rob_idx] && soc2.core.jmp_unit.imul.r_uops_1_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.imul.r_uops_1_rob_idx] : 1'b1) &&
	  (soc2.core.jmp_unit.imul.r_valids_2 ? rob_valids_2[soc2.core.jmp_unit.imul.r_uops_2_rob_idx] && soc2.core.jmp_unit.imul.r_uops_2_br_mask == rob_branch_masks_2[soc2.core.jmp_unit.imul.r_uops_2_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_0.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_1.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_2.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_3.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_4.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_5.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_6.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_7.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_8.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_9.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_10.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_11.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_12.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_13.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_14.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fp_issue_unit.slots_15.io_valid /*&& !(soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx] && soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.queue.valids_0 /*&& !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.queue.valids_1 /*&& !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.queue.valids_2 /*&& !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.queue.valids_3 /*&& !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.queue.valids_4 /*&& !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.queue.valids_5 /*&& !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.queue.valids_6 /*&& !(soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0 ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1 ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2 ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_val ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_val ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_0 && !(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_stq_idx]) ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_1 && !(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_stq_idx]) ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_2 && !(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_stq_idx]) ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_3 && !(soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_stq_idx]) ? rob_valids_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx] && soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fregister_read.exe_reg_valids_0 /*&& !(soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx] && soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx] : 1'b1) &&
	  (soc2.core.fp_pipeline.fregister_read.rrd_valids_0_REG /*&& !(soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_stq_idx]) */? rob_valids_2[soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx] && soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_br_mask == rob_branch_masks_2[soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_0.io_valid /*&& !(soc2.core.int_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_0.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_0.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_0.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_0.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_1.io_valid /*&& !(soc2.core.int_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_1.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_1.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_1.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_1.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_2.io_valid /*&& !(soc2.core.int_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_2.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_2.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_2.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_2.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_3.io_valid /*&& !(soc2.core.int_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_3.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_3.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_3.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_3.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_4.io_valid /*&& !(soc2.core.int_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_4.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_4.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_4.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_4.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_5.io_valid /*&& !(soc2.core.int_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_5.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_5.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_5.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_5.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_6.io_valid /*&& !(soc2.core.int_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_6.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_6.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_6.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_6.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_7.io_valid /*&& !(soc2.core.int_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_7.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_7.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_7.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_7.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_8.io_valid /*&& !(soc2.core.int_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_8.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_8.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_8.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_8.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_9.io_valid /*&& !(soc2.core.int_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_9.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_9.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_9.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_9.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_10.io_valid /*&& !(soc2.core.int_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_10.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_10.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_10.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_10.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_11.io_valid /*&& !(soc2.core.int_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_11.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_11.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_11.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_11.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_12.io_valid /*&& !(soc2.core.int_issue_unit.slots_12.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_12.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_12.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_12.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_12.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_13.io_valid /*&& !(soc2.core.int_issue_unit.slots_13.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_13.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_13.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_13.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_13.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_14.io_valid /*&& !(soc2.core.int_issue_unit.slots_14.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_14.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_14.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_14.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_14.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_15.io_valid /*&& !(soc2.core.int_issue_unit.slots_15.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_15.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_15.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_15.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_15.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_16.io_valid /*&& !(soc2.core.int_issue_unit.slots_16.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_16.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_16.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_16.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_16.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_17.io_valid /*&& !(soc2.core.int_issue_unit.slots_17.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_17.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_17.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_17.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_17.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_18.io_valid /*&& !(soc2.core.int_issue_unit.slots_18.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_18.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_18.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_18.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_18.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.int_issue_unit.slots_19.io_valid /*&& !(soc2.core.int_issue_unit.slots_19.slot_uop_uses_stq && stq_committed_2[soc2.core.int_issue_unit.slots_19.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.int_issue_unit.slots_19.slot_uop_rob_idx] && soc2.core.int_issue_unit.slots_19.slot_uop_br_mask == rob_branch_masks_2[soc2.core.int_issue_unit.slots_19.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_0.io_valid /*&& !(soc2.core.mem_issue_unit.slots_0.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_0.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_0.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_0.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_0.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_1.io_valid /*&& !(soc2.core.mem_issue_unit.slots_1.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_1.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_1.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_1.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_1.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_2.io_valid /*&& !(soc2.core.mem_issue_unit.slots_2.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_2.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_2.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_2.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_2.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_3.io_valid /*&& !(soc2.core.mem_issue_unit.slots_3.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_3.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_3.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_3.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_3.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_4.io_valid /*&& !(soc2.core.mem_issue_unit.slots_4.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_4.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_4.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_4.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_4.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_5.io_valid /*&& !(soc2.core.mem_issue_unit.slots_5.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_5.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_5.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_5.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_5.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_6.io_valid /*&& !(soc2.core.mem_issue_unit.slots_6.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_6.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_6.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_6.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_6.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_7.io_valid /*&& !(soc2.core.mem_issue_unit.slots_7.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_7.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_7.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_7.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_7.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_8.io_valid /*&& !(soc2.core.mem_issue_unit.slots_8.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_8.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_8.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_8.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_8.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_9.io_valid /*&& !(soc2.core.mem_issue_unit.slots_9.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_9.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_9.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_9.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_9.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_10.io_valid /*&& !(soc2.core.mem_issue_unit.slots_10.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_10.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_10.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_10.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_10.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.core.mem_issue_unit.slots_11.io_valid /*&& !(soc2.core.mem_issue_unit.slots_11.slot_uop_uses_stq && stq_committed_2[soc2.core.mem_issue_unit.slots_11.slot_uop_stq_idx]) */? rob_valids_2[soc2.core.mem_issue_unit.slots_11.slot_uop_rob_idx] && soc2.core.mem_issue_unit.slots_11.slot_uop_br_mask == rob_branch_masks_2[soc2.core.mem_issue_unit.slots_11.slot_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_0_valid ? rob_valids_2[soc2.lsu.ldq_0_bits_uop_rob_idx] && soc2.lsu.ldq_0_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_0_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_1_valid ? rob_valids_2[soc2.lsu.ldq_1_bits_uop_rob_idx] && soc2.lsu.ldq_1_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_1_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_2_valid ? rob_valids_2[soc2.lsu.ldq_2_bits_uop_rob_idx] && soc2.lsu.ldq_2_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_2_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_3_valid ? rob_valids_2[soc2.lsu.ldq_3_bits_uop_rob_idx] && soc2.lsu.ldq_3_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_3_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_4_valid ? rob_valids_2[soc2.lsu.ldq_4_bits_uop_rob_idx] && soc2.lsu.ldq_4_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_4_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_5_valid ? rob_valids_2[soc2.lsu.ldq_5_bits_uop_rob_idx] && soc2.lsu.ldq_5_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_5_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_6_valid ? rob_valids_2[soc2.lsu.ldq_6_bits_uop_rob_idx] && soc2.lsu.ldq_6_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_6_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_7_valid ? rob_valids_2[soc2.lsu.ldq_7_bits_uop_rob_idx] && soc2.lsu.ldq_7_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_7_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_8_valid ? rob_valids_2[soc2.lsu.ldq_8_bits_uop_rob_idx] && soc2.lsu.ldq_8_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_8_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_9_valid ? rob_valids_2[soc2.lsu.ldq_9_bits_uop_rob_idx] && soc2.lsu.ldq_9_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_9_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_10_valid ? rob_valids_2[soc2.lsu.ldq_10_bits_uop_rob_idx] && soc2.lsu.ldq_10_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_10_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_11_valid ? rob_valids_2[soc2.lsu.ldq_11_bits_uop_rob_idx] && soc2.lsu.ldq_11_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_11_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_12_valid ? rob_valids_2[soc2.lsu.ldq_12_bits_uop_rob_idx] && soc2.lsu.ldq_12_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_12_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_13_valid ? rob_valids_2[soc2.lsu.ldq_13_bits_uop_rob_idx] && soc2.lsu.ldq_13_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_13_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_14_valid ? rob_valids_2[soc2.lsu.ldq_14_bits_uop_rob_idx] && soc2.lsu.ldq_14_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_14_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_15_valid ? rob_valids_2[soc2.lsu.ldq_15_bits_uop_rob_idx] && soc2.lsu.ldq_15_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.ldq_15_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.fired_sfence_0 ? rob_valids_2[soc2.lsu.mem_incoming_uop_0_rob_idx] && soc2.lsu.mem_incoming_uop_0_br_mask == rob_branch_masks_2[soc2.lsu.mem_incoming_uop_0_rob_idx] : 1'b1) &&
	  ((soc2.lsu.fired_stad_incoming_REG || soc2.lsu.fired_sta_incoming_REG || soc2.lsu.fired_std_incoming_REG) /*&& !stq_committed_2[soc2.lsu.mem_stq_incoming_e_0_bits_uop_stq_idx] */? rob_valids_2[soc2.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx] && soc2.lsu.mem_stq_incoming_e_0_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.fired_sta_retry_REG /*&& !stq_committed_2[soc2.lsu.mem_stq_retry_e_bits_uop_stq_idx] */? rob_valids_2[soc2.lsu.mem_stq_retry_e_bits_uop_rob_idx] && soc2.lsu.mem_stq_retry_e_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.mem_stq_retry_e_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.mem_xcpt_valids_0 /*&& !(soc2.lsu.mem_xcpt_uops_0_uses_stq && stq_committed_2[soc2.lsu.mem_xcpt_uops_0_stq_idx]) */? rob_valids_2[soc2.lsu.mem_xcpt_uops_0_rob_idx] && soc2.lsu.mem_xcpt_uops_0_br_mask == rob_branch_masks_2[soc2.lsu.mem_xcpt_uops_0_rob_idx] : 1'b1) &&
	  (soc2.lsu.fired_stdf_incoming /*&& !stq_committed_2[soc2.lsu.mem_stdf_uop_stq_idx] */? rob_valids_2[soc2.lsu.mem_stdf_uop_rob_idx] && soc2.lsu.mem_stdf_uop_br_mask == rob_branch_masks_2[soc2.lsu.mem_stdf_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stdf_clr_bsy_valid ? rob_valids_2[soc2.lsu.stdf_clr_bsy_rob_idx] && soc2.lsu.stdf_clr_bsy_brmask == rob_branch_masks_2[soc2.lsu.stdf_clr_bsy_rob_idx] : 1'b1) &&
	  //stores do not have to be checked after they are committed (their ROB entry can be used for another uop then)
	  (soc2.lsu.stq_0_valid && !soc2.lsu.stq_0_bits_committed ? rob_valids_2[soc2.lsu.stq_0_bits_uop_rob_idx] && soc2.lsu.stq_0_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_0_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_1_valid && !soc2.lsu.stq_1_bits_committed ? rob_valids_2[soc2.lsu.stq_1_bits_uop_rob_idx] && soc2.lsu.stq_1_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_1_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_2_valid && !soc2.lsu.stq_2_bits_committed ? rob_valids_2[soc2.lsu.stq_2_bits_uop_rob_idx] && soc2.lsu.stq_2_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_2_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_3_valid && !soc2.lsu.stq_3_bits_committed ? rob_valids_2[soc2.lsu.stq_3_bits_uop_rob_idx] && soc2.lsu.stq_3_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_3_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_4_valid && !soc2.lsu.stq_4_bits_committed ? rob_valids_2[soc2.lsu.stq_4_bits_uop_rob_idx] && soc2.lsu.stq_4_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_4_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_5_valid && !soc2.lsu.stq_5_bits_committed ? rob_valids_2[soc2.lsu.stq_5_bits_uop_rob_idx] && soc2.lsu.stq_5_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_5_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_6_valid && !soc2.lsu.stq_6_bits_committed ? rob_valids_2[soc2.lsu.stq_6_bits_uop_rob_idx] && soc2.lsu.stq_6_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_6_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_7_valid && !soc2.lsu.stq_7_bits_committed ? rob_valids_2[soc2.lsu.stq_7_bits_uop_rob_idx] && soc2.lsu.stq_7_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_7_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_8_valid && !soc2.lsu.stq_8_bits_committed ? rob_valids_2[soc2.lsu.stq_8_bits_uop_rob_idx] && soc2.lsu.stq_8_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_8_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_9_valid && !soc2.lsu.stq_9_bits_committed ? rob_valids_2[soc2.lsu.stq_9_bits_uop_rob_idx] && soc2.lsu.stq_9_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_9_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_10_valid && !soc2.lsu.stq_10_bits_committed ? rob_valids_2[soc2.lsu.stq_10_bits_uop_rob_idx] && soc2.lsu.stq_10_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_10_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_11_valid && !soc2.lsu.stq_11_bits_committed ? rob_valids_2[soc2.lsu.stq_11_bits_uop_rob_idx] && soc2.lsu.stq_11_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_11_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_12_valid && !soc2.lsu.stq_12_bits_committed ? rob_valids_2[soc2.lsu.stq_12_bits_uop_rob_idx] && soc2.lsu.stq_12_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_12_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_13_valid && !soc2.lsu.stq_13_bits_committed ? rob_valids_2[soc2.lsu.stq_13_bits_uop_rob_idx] && soc2.lsu.stq_13_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_13_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_14_valid && !soc2.lsu.stq_14_bits_committed ? rob_valids_2[soc2.lsu.stq_14_bits_uop_rob_idx] && soc2.lsu.stq_14_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_14_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.stq_15_valid && !soc2.lsu.stq_15_bits_committed ? rob_valids_2[soc2.lsu.stq_15_bits_uop_rob_idx] && soc2.lsu.stq_15_bits_uop_br_mask == rob_branch_masks_2[soc2.lsu.stq_15_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.clr_bsy_valid_0 ? rob_valids_2[soc2.lsu.clr_bsy_rob_idx_0] && soc2.lsu.clr_bsy_brmask_0 == rob_branch_masks_2[soc2.lsu.clr_bsy_rob_idx_0] : 1'b1) &&
	  (soc2.lsu.r_xcpt_valid ? rob_valids_2[soc2.lsu.r_xcpt_uop_rob_idx] && soc2.lsu.r_xcpt_uop_br_mask == rob_branch_masks_2[soc2.lsu.r_xcpt_uop_rob_idx] : 1'b1) &&

	  (soc2.dcache.mshrs.respq.valids_0
	  ? (
	    (soc2.dcache.mshrs.respq.uops_0_uses_ldq ? rob_valids_2[ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_0_ldq_idx]] && soc2.dcache.mshrs.respq.uops_0_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_0_ldq_idx]] : 1'b1) &&
	    (soc2.dcache.mshrs.respq.uops_0_uses_stq && !stq_committed_2[soc2.dcache.mshrs.respq.uops_0_stq_idx] ? rob_valids_2[stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_0_stq_idx]] && soc2.dcache.mshrs.respq.uops_0_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_0_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.respq.valids_1
	  ? (
	    (soc2.dcache.mshrs.respq.uops_1_uses_ldq ? rob_valids_2[ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_1_ldq_idx]] && soc2.dcache.mshrs.respq.uops_1_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_1_ldq_idx]] : 1'b1) &&
	    (soc2.dcache.mshrs.respq.uops_1_uses_stq && !stq_committed_2[soc2.dcache.mshrs.respq.uops_1_stq_idx] ? rob_valids_2[stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_1_stq_idx]] && soc2.dcache.mshrs.respq.uops_1_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_1_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.respq.valids_2
	  ? (
	    (soc2.dcache.mshrs.respq.uops_2_uses_ldq ? rob_valids_2[ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_2_ldq_idx]] && soc2.dcache.mshrs.respq.uops_2_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_2_ldq_idx]] : 1'b1) &&
	    (soc2.dcache.mshrs.respq.uops_2_uses_stq && !stq_committed_2[soc2.dcache.mshrs.respq.uops_2_stq_idx] ? rob_valids_2[stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_2_stq_idx]] && soc2.dcache.mshrs.respq.uops_2_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_2_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.respq.valids_3
	  ? (
	    (soc2.dcache.mshrs.respq.uops_3_uses_ldq ? rob_valids_2[ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_3_ldq_idx]] && soc2.dcache.mshrs.respq.uops_3_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.respq.uops_3_ldq_idx]] : 1'b1) &&
	    (soc2.dcache.mshrs.respq.uops_3_uses_stq && !stq_committed_2[soc2.dcache.mshrs.respq.uops_3_stq_idx] ? rob_valids_2[stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_3_stq_idx]] && soc2.dcache.mshrs.respq.uops_3_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.respq.uops_3_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mmios_0.state != 2'b0
	  ? (
	    (soc2.dcache.mshrs.mmios_0.req_uop_uses_ldq ? rob_valids_2[ldq_rob_idx_2[soc2.dcache.mshrs.mmios_0.req_uop_ldq_idx]] && soc2.dcache.mshrs.mmios_0.req_uop_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mmios_0.req_uop_ldq_idx]] : 1'b1) &&
	    (soc2.dcache.mshrs.mmios_0.req_uop_uses_stq && !stq_committed_2[soc2.dcache.mshrs.mmios_0.req_uop_stq_idx] ? rob_valids_2[stq_rob_idx_2[soc2.dcache.mshrs.mmios_0.req_uop_stq_idx]] && soc2.dcache.mshrs.mmios_0.req_uop_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mmios_0.req_uop_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_0
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_0_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_0_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_0_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_1
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_1_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_1_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_1_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_2
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_2_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_2_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_2_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_3
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_3_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_3_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_3_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_4
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_4_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_4_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_4_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_5
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_5_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_5_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_5_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_6
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_6_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_6_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_6_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_7
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_7_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_7_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_7_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_8
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_8_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_8_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_8_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_9
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_9_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_9_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_9_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_10
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_10_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_10_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_10_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_11
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_11_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_11_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_11_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_12
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_12_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_12_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_12_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_13
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_13_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_13_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_13_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_14
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_14_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_14_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_14_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_15
	  ? (
	    (soc2.dcache.mshrs.mshrs_0.rpq.uops_15_uses_ldq ? soc2.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_15_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_0.rpq.uops_15_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx] ? soc2.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_0
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_0_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_0_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_0_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_1
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_1_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_1_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_1_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_2
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_2_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_2_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_2_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_3
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_3_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_3_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_3_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_4
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_4_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_4_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_4_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_5
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_5_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_5_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_5_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_6
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_6_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_6_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_6_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_7
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_7_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_7_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_7_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_8
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_8_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_8_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_8_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_9
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_9_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_9_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_9_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_10
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_10_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_10_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_10_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_11
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_11_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_11_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_11_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_12
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_12_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_12_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_12_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_13
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_13_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_13_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_13_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_14
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_14_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_14_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_14_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_15
	  ? (
	    (soc2.dcache.mshrs.mshrs_1.rpq.uops_15_uses_ldq ? soc2.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_15_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.mshrs.mshrs_1.rpq.uops_15_uses_stq && !stq_committed[soc2.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx] ? soc2.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.s1_valid_REG
	  ? (
	    (soc2.dcache.s1_req_0_uop_uses_ldq ? soc2.dcache.s1_req_0_uop_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.s1_req_0_uop_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.s1_req_0_uop_uses_stq ? soc2.dcache.s1_req_0_uop_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.s1_req_0_uop_stq_idx]] : 1'b1))
	  :
	    1'b1) &&
	  (soc2.dcache.s2_valid_REG
	  ? (
	    (soc2.dcache.s2_req_0_uop_uses_ldq ? soc2.dcache.s2_req_0_uop_br_mask == rob_branch_masks_2[ldq_rob_idx_2[soc2.dcache.s2_req_0_uop_ldq_idx]] : 1'b1) //&&
	    )//(soc2.dcache.s2_req_0_uop_uses_stq ? soc2.dcache.s2_req_0_uop_br_mask == rob_branch_masks_2[stq_rob_idx_2[soc2.dcache.s2_req_0_uop_stq_idx]] : 1'b1))
	  :
	    1'b1)
	  ;

	//check for all issue slots:
	//if the corresponding ROB entry is invalid the state of the issue slot has to be invalid too
	wire valid_issue_slots_2;
	assign valid_issue_slots_2 =
	(!rob_valids_2[soc2.core.int_issue_unit.slots_0.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_0.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_1.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_1.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_2.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_2.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_3.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_3.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_4.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_4.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_5.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_5.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_6.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_6.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_7.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_7.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_8.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_8.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_9.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_9.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_10.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_10.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_11.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_11.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_12.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_12.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_13.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_13.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_14.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_14.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_15.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_15.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_16.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_16.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_17.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_17.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_18.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_18.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.int_issue_unit.slots_19.slot_uop_rob_idx] ? soc2.core.int_issue_unit.slots_19.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_0.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_0.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_1.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_1.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_2.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_2.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_3.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_3.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_4.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_4.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_5.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_5.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_6.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_6.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_7.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_7.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_8.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_8.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_9.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_9.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_10.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_10.state == 2'b0 : 1'b1) &&
	(!rob_valids_2[soc2.core.mem_issue_unit.slots_11.slot_uop_rob_idx] ? soc2.core.mem_issue_unit.slots_11.state == 2'b0 : 1'b1);

	//check for the branch misprediction:
	//if the prediction is valid the corresponding ROB entry must be valid too
	wire valid_mispred_idx_2;
	assign valid_mispred_idx_2 =
	(soc2.core.brinfos_0_valid ? rob_valids_2[soc2.core.brinfos_0_uop_rob_idx] : 1'b1) &&
	(soc2.core.brinfos_1_valid ? rob_valids_2[soc2.core.brinfos_1_uop_rob_idx] : 1'b1);

	//check for iregister read buffers:
	//if the buffer is valid the corresponding ROB entry must be valid too
	wire valid_iregister_read_2;
	assign valid_iregister_read_2 =
	(soc2.core.iregister_read.exe_reg_valids_1 ? rob_valids_2[soc2.core.iregister_read.exe_reg_uops_1_rob_idx] : 1'b1) &&
	(soc2.core.iregister_read.exe_reg_valids_2 ? rob_valids_2[soc2.core.iregister_read.exe_reg_uops_2_rob_idx] : 1'b1) &&
	(soc2.core.iregister_read.rrd_valids_1_REG ? rob_valids_2[soc2.core.iregister_read.rrd_uops_1_REG_rob_idx] : 1'b1) &&
	(soc2.core.iregister_read.rrd_valids_2_REG ? rob_valids_2[soc2.core.iregister_read.rrd_uops_2_REG_rob_idx] : 1'b1);

	//instruction at head must be non-speculative (br_mask == 0) if it is valid
	wire no_speculative_head_2;
	assign no_speculative_head_2 =
	  rob_valids_2[soc2.core.rob.io_rob_head_idx]? (rob_branch_masks_2[soc2.core.rob.io_rob_head_idx] == 12'b0) : 1'b1;

	//ensure that valid entries are not overwritten
	wire prevent_overwriting_valid_entries_2;
	assign prevent_overwriting_valid_entries_2 = 
		(soc2.core.rob.io_enq_valids_0 ? !rob_valids_2[{soc2.core.rob.rob_tail,1'b0}] : 1'b1) &&
		(soc2.core.rob.io_enq_valids_1 ? !rob_valids_2[{soc2.core.rob.rob_tail,1'b1}] : 1'b1);
		
	//ROB is never full and empty
	wire full_empty_logic_2;
	assign full_empty_logic_2 = !(soc2.core.rob.full && soc2.core.rob.empty);

	//ROB is empty equals head == tail and all valid bits are 0
	wire empty_logic_2;
	assign empty_logic_2 =
	  ((soc2.core.rob.rob_head == soc2.core.rob.rob_tail) && ((rob_valids_2[0] | rob_valids_2[1] | rob_valids_2[2] | rob_valids_2[3] | rob_valids_2[4] | rob_valids_2[5] | rob_valids_2[6] | rob_valids_2[7] | rob_valids_2[8] | rob_valids_2[9] |
	    rob_valids_2[10] | rob_valids_2[11] | rob_valids_2[12] | rob_valids_2[13] | rob_valids_2[14] | rob_valids_2[15] | rob_valids_2[16] | rob_valids_2[17] | rob_valids_2[18] | rob_valids_2[19] | 
	    rob_valids_2[20] | rob_valids_2[21] | rob_valids_2[22] | rob_valids_2[23] | rob_valids_2[24] | rob_valids_2[25] | rob_valids_2[26] | rob_valids_2[27] | rob_valids_2[28] | rob_valids_2[29] | 
	    rob_valids_2[30] | rob_valids_2[31] | rob_valids_2[32] | rob_valids_2[33] | rob_valids_2[34] | rob_valids_2[35] | rob_valids_2[36] | rob_valids_2[37] | rob_valids_2[38] | rob_valids_2[39] | 
	    rob_valids_2[40] | rob_valids_2[41] | rob_valids_2[42] | rob_valids_2[43] | rob_valids_2[44] | rob_valids_2[45] | rob_valids_2[46] | rob_valids_2[47] | rob_valids_2[48] | rob_valids_2[49] | 
	    rob_valids_2[50] | rob_valids_2[51] | rob_valids_2[52] | rob_valids_2[53] | rob_valids_2[54] | rob_valids_2[55] | rob_valids_2[56] | rob_valids_2[57] | rob_valids_2[58] | rob_valids_2[59] | 
	    rob_valids_2[60] | rob_valids_2[61] | rob_valids_2[62] | rob_valids_2[63]) == 1'b0)) == soc2.core.rob.empty;
	    
	//ROB is full equals head == tail and either one of the entrys at tail is valid or tail_lsb is not set, else rob_state is rollback
	wire full_logic_2;
	assign full_logic_2 = (soc2.core.rob.rob_head == soc2.core.rob.rob_tail && soc2.core.rob.maybe_full) == soc2.core.rob.full;
	  
	//Create array for load queue valid bits
	wire ldq_valids_2 [15:0];
	assign ldq_valids_2[0] = soc2.lsu.ldq_0_valid;
	assign ldq_valids_2[1] = soc2.lsu.ldq_1_valid;
	assign ldq_valids_2[2] = soc2.lsu.ldq_2_valid;
	assign ldq_valids_2[3] = soc2.lsu.ldq_3_valid;
	assign ldq_valids_2[4] = soc2.lsu.ldq_4_valid;
	assign ldq_valids_2[5] = soc2.lsu.ldq_5_valid;
	assign ldq_valids_2[6] = soc2.lsu.ldq_6_valid;
	assign ldq_valids_2[7] = soc2.lsu.ldq_7_valid;
	assign ldq_valids_2[8] = soc2.lsu.ldq_8_valid;
	assign ldq_valids_2[9] = soc2.lsu.ldq_9_valid;
	assign ldq_valids_2[10] = soc2.lsu.ldq_10_valid;
	assign ldq_valids_2[11] = soc2.lsu.ldq_11_valid;
	assign ldq_valids_2[12] = soc2.lsu.ldq_12_valid;
	assign ldq_valids_2[13] = soc2.lsu.ldq_13_valid;
	assign ldq_valids_2[14] = soc2.lsu.ldq_14_valid;
	assign ldq_valids_2[15] = soc2.lsu.ldq_15_valid;
	  
	wire lcam_ldq_idx_valid_2;
	assign lcam_ldq_idx_valid_2 = 
	//if a load got fired, its ldq entry has to be valid
	(soc2.lsu.fired_load_incoming_REG || soc2.lsu.fired_load_retry_REG || soc2.lsu.fired_load_wakeup_REG) && !soc2.lsu.REG_1 ? ldq_valids_2[soc2.lsu.lcam_ldq_idx_0] : 1'b1;
	
	//Create array for load queue valid bits
	wire stq_valids_2 [15:0];
	assign stq_valids_2[0] = soc2.lsu.stq_0_valid;
	assign stq_valids_2[1] = soc2.lsu.stq_1_valid;
	assign stq_valids_2[2] = soc2.lsu.stq_2_valid;
	assign stq_valids_2[3] = soc2.lsu.stq_3_valid;
	assign stq_valids_2[4] = soc2.lsu.stq_4_valid;
	assign stq_valids_2[5] = soc2.lsu.stq_5_valid;
	assign stq_valids_2[6] = soc2.lsu.stq_6_valid;
	assign stq_valids_2[7] = soc2.lsu.stq_7_valid;
	assign stq_valids_2[8] = soc2.lsu.stq_8_valid;
	assign stq_valids_2[9] = soc2.lsu.stq_9_valid;
	assign stq_valids_2[10] = soc2.lsu.stq_10_valid;
	assign stq_valids_2[11] = soc2.lsu.stq_11_valid;
	assign stq_valids_2[12] = soc2.lsu.stq_12_valid;
	assign stq_valids_2[13] = soc2.lsu.stq_13_valid;
	assign stq_valids_2[14] = soc2.lsu.stq_14_valid;
	assign stq_valids_2[15] = soc2.lsu.stq_15_valid;

	wire lcam_stq_idx_valid_2;
	assign lcam_stq_idx_valid_2 = 
	//if a load got fired, its stq entry has to be valid
	(soc2.lsu.fired_sta_incoming_REG || soc2.lsu.fired_stad_incoming_REG || soc2.lsu.fired_sta_retry_REG) && !soc2.lsu.REG_1 ? stq_valids_2[soc2.lsu.lcam_stq_idx_0] : 1'b1;
	  
	  
	wire ldq_consistent_rob_idx_2;
	assign ldq_consistent_rob_idx_2 =
	  (ldq_valids_2[soc2.lsu.ldq_head])
	  ?
	    (ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 0) % 16], soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx) ? 1'b1 : (soc2.core.rob.full && (soc2.core.rob.io_rob_head_idx == soc2.core.rob.io_rob_tail_idx))) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 1) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 0) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 1) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 2) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 1) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 2) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 3) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 2) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 3) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 4) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 3) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 4) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 5) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 4) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 5) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 6) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 5) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 6) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 7) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 6) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 7) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 8) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 7) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 8) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 9) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 8) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 9) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 10) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 9) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 10) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 11) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 10) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 11) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 12) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 11) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 12) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 13) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 12) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 13) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 14) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 13) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 14) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (ldq_valids_2[(soc2.lsu.ldq_head + 15) % 16] ? ROBisOlder(ldq_rob_idx_2[(soc2.lsu.ldq_head + 14) % 16], ldq_rob_idx_2[(soc2.lsu.ldq_head + 15) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1)
	  :
	  	1'b1;

	wire stq_consistent_rob_idx_2;
	assign stq_consistent_rob_idx_2 =
	  stq_valids_2[soc2.lsu.stq_head]
		  ?
	    (ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 0) % 16], soc2.core.rob.io_rob_tail_idx, soc2.core.rob.io_rob_head_idx) ? 1'b1 : (stq_committed_2[(soc2.lsu.stq_head + 0) % 16]) || (soc2.core.rob.full && (soc2.core.rob.io_rob_head_idx == soc2.core.rob.io_rob_tail_idx))) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 1) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 1) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 0) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 0) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 1) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 2) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 2) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 1) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 1) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 2) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 3) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 3) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 2) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 2) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 3) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 4) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 4) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 3) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 3) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 4) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 5) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 5) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 4) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 4) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 5) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 6) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 6) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 5) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 5) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 6) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 7) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 7) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 6) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 6) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 7) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 8) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 8) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 7) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 7) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 8) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 9) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 9) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 8) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 8) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 9) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 10) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 10) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 9) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 9) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 10) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 11) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 11) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 10) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 10) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 11) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 12) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 12) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 11) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 11) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 12) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 13) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 13) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 12) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 12) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 13) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 14) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 14) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 13) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 13) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 14) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	    (stq_valids_2[(soc2.lsu.stq_head + 15) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 15) % 16] && !stq_committed_2[(soc2.lsu.stq_head + 14) % 16] ? ROBisOlder(stq_rob_idx_2[(soc2.lsu.stq_head + 14) % 16], stq_rob_idx_2[(soc2.lsu.stq_head + 15) % 16], soc2.core.rob.io_rob_head_idx) : 1'b1)
	  :
	  	1'b1;  
	  
	wire consistent_stq_committed_2;
	assign consistent_stq_committed_2 =
	(soc2.lsu.stq_0_bits_committed ? soc2.lsu.stq_0_valid : 1'b1) &&
	(soc2.lsu.stq_1_bits_committed ? soc2.lsu.stq_1_valid : 1'b1) &&
	(soc2.lsu.stq_2_bits_committed ? soc2.lsu.stq_2_valid : 1'b1) &&
	(soc2.lsu.stq_3_bits_committed ? soc2.lsu.stq_3_valid : 1'b1) &&
	(soc2.lsu.stq_4_bits_committed ? soc2.lsu.stq_4_valid : 1'b1) &&
	(soc2.lsu.stq_5_bits_committed ? soc2.lsu.stq_5_valid : 1'b1) &&
	(soc2.lsu.stq_6_bits_committed ? soc2.lsu.stq_6_valid : 1'b1) &&
	(soc2.lsu.stq_7_bits_committed ? soc2.lsu.stq_7_valid : 1'b1) &&
	(soc2.lsu.stq_8_bits_committed ? soc2.lsu.stq_8_valid : 1'b1) &&
	(soc2.lsu.stq_9_bits_committed ? soc2.lsu.stq_9_valid : 1'b1) &&
	(soc2.lsu.stq_10_bits_committed ? soc2.lsu.stq_10_valid : 1'b1) &&
	(soc2.lsu.stq_11_bits_committed ? soc2.lsu.stq_11_valid : 1'b1) &&
	(soc2.lsu.stq_12_bits_committed ? soc2.lsu.stq_12_valid : 1'b1) &&
	(soc2.lsu.stq_13_bits_committed ? soc2.lsu.stq_13_valid : 1'b1) &&
	(soc2.lsu.stq_14_bits_committed ? soc2.lsu.stq_14_valid : 1'b1) &&
	(soc2.lsu.stq_15_bits_committed ? soc2.lsu.stq_15_valid : 1'b1);
	
	wire committed_stores_not_speculative_2;
	assign committed_stores_not_speculative_2 =
	  (soc2.lsu.stq_0_bits_committed ? soc2.lsu.stq_0_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_1_bits_committed ? soc2.lsu.stq_1_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_2_bits_committed ? soc2.lsu.stq_2_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_3_bits_committed ? soc2.lsu.stq_3_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_4_bits_committed ? soc2.lsu.stq_4_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_5_bits_committed ? soc2.lsu.stq_5_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_6_bits_committed ? soc2.lsu.stq_6_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_7_bits_committed ? soc2.lsu.stq_7_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_8_bits_committed ? soc2.lsu.stq_8_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_9_bits_committed ? soc2.lsu.stq_9_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_10_bits_committed ? soc2.lsu.stq_10_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_11_bits_committed ? soc2.lsu.stq_11_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_12_bits_committed ? soc2.lsu.stq_12_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_13_bits_committed ? soc2.lsu.stq_13_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_14_bits_committed ? soc2.lsu.stq_14_bits_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.lsu.stq_15_bits_committed ? soc2.lsu.stq_15_bits_uop_br_mask == 12'b0 : 1'b1);

	wire ldq_rob_valid_consistency_2;
	assign ldq_rob_valid_consistency_2 =
	  (soc2.lsu.ldq_0_valid ? rob_valids_2[soc2.lsu.ldq_0_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_1_valid ? rob_valids_2[soc2.lsu.ldq_1_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_2_valid ? rob_valids_2[soc2.lsu.ldq_2_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_3_valid ? rob_valids_2[soc2.lsu.ldq_3_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_4_valid ? rob_valids_2[soc2.lsu.ldq_4_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_5_valid ? rob_valids_2[soc2.lsu.ldq_5_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_6_valid ? rob_valids_2[soc2.lsu.ldq_6_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_7_valid ? rob_valids_2[soc2.lsu.ldq_7_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_8_valid ? rob_valids_2[soc2.lsu.ldq_8_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_9_valid ? rob_valids_2[soc2.lsu.ldq_9_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_10_valid ? rob_valids_2[soc2.lsu.ldq_10_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_11_valid ? rob_valids_2[soc2.lsu.ldq_11_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_12_valid ? rob_valids_2[soc2.lsu.ldq_12_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_13_valid ? rob_valids_2[soc2.lsu.ldq_13_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_14_valid ? rob_valids_2[soc2.lsu.ldq_14_bits_uop_rob_idx] : 1'b1) &&
	  (soc2.lsu.ldq_15_valid ? rob_valids_2[soc2.lsu.ldq_15_bits_uop_rob_idx] : 1'b1);

	wire speculative_store_rpq_2;
	assign speculative_store_rpq_2 =
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_0 && soc2.dcache.mshrs.mshrs_0.rpq.uops_0_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_0_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_1 && soc2.dcache.mshrs.mshrs_0.rpq.uops_1_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_1_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_2 && soc2.dcache.mshrs.mshrs_0.rpq.uops_2_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_2_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_3 && soc2.dcache.mshrs.mshrs_0.rpq.uops_3_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_3_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_4 && soc2.dcache.mshrs.mshrs_0.rpq.uops_4_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_4_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_5 && soc2.dcache.mshrs.mshrs_0.rpq.uops_5_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_5_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_6 && soc2.dcache.mshrs.mshrs_0.rpq.uops_6_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_6_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_7 && soc2.dcache.mshrs.mshrs_0.rpq.uops_7_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_7_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_8 && soc2.dcache.mshrs.mshrs_0.rpq.uops_8_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_8_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_9 && soc2.dcache.mshrs.mshrs_0.rpq.uops_9_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_9_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_10 && soc2.dcache.mshrs.mshrs_0.rpq.uops_10_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_10_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_11 && soc2.dcache.mshrs.mshrs_0.rpq.uops_11_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_11_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_12 && soc2.dcache.mshrs.mshrs_0.rpq.uops_12_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_12_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_13 && soc2.dcache.mshrs.mshrs_0.rpq.uops_13_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_13_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_14 && soc2.dcache.mshrs.mshrs_0.rpq.uops_14_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_14_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_0.rpq.valids_15 && soc2.dcache.mshrs.mshrs_0.rpq.uops_15_uses_stq && (soc2.dcache.mshrs.mshrs_0.rpq.uops_15_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_0 && soc2.dcache.mshrs.mshrs_1.rpq.uops_0_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_0_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_1 && soc2.dcache.mshrs.mshrs_1.rpq.uops_1_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_1_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_2 && soc2.dcache.mshrs.mshrs_1.rpq.uops_2_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_2_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_3 && soc2.dcache.mshrs.mshrs_1.rpq.uops_3_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_3_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_4 && soc2.dcache.mshrs.mshrs_1.rpq.uops_4_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_4_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_5 && soc2.dcache.mshrs.mshrs_1.rpq.uops_5_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_5_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_6 && soc2.dcache.mshrs.mshrs_1.rpq.uops_6_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_6_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_7 && soc2.dcache.mshrs.mshrs_1.rpq.uops_7_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_7_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_8 && soc2.dcache.mshrs.mshrs_1.rpq.uops_8_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_8_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_9 && soc2.dcache.mshrs.mshrs_1.rpq.uops_9_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_9_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_10 && soc2.dcache.mshrs.mshrs_1.rpq.uops_10_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_10_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_11 && soc2.dcache.mshrs.mshrs_1.rpq.uops_11_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_11_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_12 && soc2.dcache.mshrs.mshrs_1.rpq.uops_12_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_12_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_13 && soc2.dcache.mshrs.mshrs_1.rpq.uops_13_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_13_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_14 && soc2.dcache.mshrs.mshrs_1.rpq.uops_14_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_14_br_mask != 12'b0)) ||
	  (soc2.dcache.mshrs.mshrs_1.rpq.valids_15 && soc2.dcache.mshrs.mshrs_1.rpq.uops_15_uses_stq && (soc2.dcache.mshrs.mshrs_1.rpq.uops_15_br_mask != 12'b0));
	  
	wire speculative_store_s1_s2_2;
	assign speculative_store_s1_s2_2 =
	  (soc2.dcache.s1_valid_REG && soc2.dcache.s1_req_0_uop_uses_stq ? soc2.dcache.s1_req_0_uop_br_mask == 12'b0 : 1'b1) &&
	  (soc2.dcache.s2_valid_REG && soc2.dcache.s2_req_0_uop_uses_stq ? soc2.dcache.s2_req_0_uop_br_mask == 12'b0 : 1'b1);
	  
	wire fpiu_BranchKillableQueue_1_not_committed_2;
	assign fpiu_BranchKillableQueue_1_not_committed_2 =
	  (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0 ? !(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_stq_idx]) : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1 ? !(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_stq_idx]) : 1'b1) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2 ? !(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_uses_stq && stq_committed_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_stq_idx]) : 1'b1);

	wire fdivsqrt_valid_consistency_2;
	assign fdivsqrt_valid_consistency_2 = soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.io_outValid_div || soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.io_outValid_sqrt ? soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val : 1'b1;

	wire div_state_2;
	assign div_state_2 = !soc2.core.reset ? (soc2.core.csr_exe_unit.div.div.state == 3'h0) || (soc2.core.csr_exe_unit.div.div.state == 3'h3) || (soc2.core.csr_exe_unit.div.div.state == 3'h7) : 1'b1;

	wire uncom_branch_resolution;
	assign uncom_branch_resolution =
        (mispred_happened_1 == 1'b0) && (mispred_happened_2 == 1'b0) ?
        ((soc1.core.brinfos_0_valid == 1'b1) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.brinfos_0_uop_rob_idx) == 1'b1) && (soc1.core.brinfos_0_uop_rob_idx == soc2.core.brinfos_0_uop_rob_idx) ?
            soc1.core.brinfos_0_mispredict == soc2.core.brinfos_0_mispredict : 1'b1) &&
        ((soc1.core.brinfos_1_valid == 1'b1) && (isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.brinfos_1_uop_rob_idx) == 1'b1) && (soc1.core.brinfos_1_uop_rob_idx == soc2.core.brinfos_1_uop_rob_idx) ?
            soc1.core.brinfos_1_mispredict == soc2.core.brinfos_1_mispredict : 1'b1)
        :
        1'b1;
        
	wire ldq_entries_not_using_stq_2;
	assign ldq_entries_not_using_stq_2 = 
	  !soc2.lsu.ldq_0_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_1_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_2_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_3_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_4_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_5_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_6_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_7_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_8_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_9_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_10_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_11_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_12_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_13_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_14_bits_uop_uses_stq &&
	  !soc2.lsu.ldq_15_bits_uop_uses_stq;

	wire stq_entries_not_using_ldq_2;
	assign stq_entries_not_using_ldq_2 = 
	  !soc2.lsu.stq_0_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_1_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_2_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_3_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_4_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_5_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_6_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_7_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_8_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_9_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_10_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_11_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_12_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_13_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_14_bits_uop_uses_ldq &&
	  !soc2.lsu.stq_15_bits_uop_uses_ldq;
        
	wire BranchKillableQueue_empty_2;
	assign BranchKillableQueue_empty_2 =
	soc2.core.b2_mispredict ||
	(soc2.core.jmp_unit.queue.io_empty ==
	(!soc2.core.jmp_unit.queue.valids_0 &&
	!soc2.core.jmp_unit.queue.valids_1 &&
	!soc2.core.jmp_unit.queue.valids_2 &&
	!soc2.core.jmp_unit.queue.valids_3 &&
	!soc2.core.jmp_unit.queue.valids_4)) &&

	(soc2.core.fp_pipeline.fpiu_unit.queue.io_empty ==
	(!soc2.core.fp_pipeline.fpiu_unit.queue.valids_0 &&
	!soc2.core.fp_pipeline.fpiu_unit.queue.valids_1 &&
	!soc2.core.fp_pipeline.fpiu_unit.queue.valids_2 &&
	!soc2.core.fp_pipeline.fpiu_unit.queue.valids_3 &&
	!soc2.core.fp_pipeline.fpiu_unit.queue.valids_4 &&
	!soc2.core.fp_pipeline.fpiu_unit.queue.valids_5 &&
	!soc2.core.fp_pipeline.fpiu_unit.queue.valids_6)) &&

	(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.io_empty ==
	(!soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0 &&
	!soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1 &&
	!soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2)) &&

	(
	  (soc2.core.jmp_unit.queue.value == 3'h0 && soc2.core.jmp_unit.queue.valids_0) ||
	  (soc2.core.jmp_unit.queue.value == 3'h1 && soc2.core.jmp_unit.queue.valids_1) ||
	  (soc2.core.jmp_unit.queue.value == 3'h2 && soc2.core.jmp_unit.queue.valids_2) ||
	  (soc2.core.jmp_unit.queue.value == 3'h3 && soc2.core.jmp_unit.queue.valids_3) ||
	  (soc2.core.jmp_unit.queue.value == 3'h4 && soc2.core.jmp_unit.queue.valids_4)
	  ?
	  !soc2.core.jmp_unit.queue.do_enq
	  :
	  1'b1
	) &&
	(
	  (soc2.core.fp_pipeline.fpiu_unit.queue.value == 3'h0 && soc2.core.fp_pipeline.fpiu_unit.queue.valids_0) ||
	  (soc2.core.fp_pipeline.fpiu_unit.queue.value == 3'h1 && soc2.core.fp_pipeline.fpiu_unit.queue.valids_1) ||
	  (soc2.core.fp_pipeline.fpiu_unit.queue.value == 3'h2 && soc2.core.fp_pipeline.fpiu_unit.queue.valids_2) ||
	  (soc2.core.fp_pipeline.fpiu_unit.queue.value == 3'h3 && soc2.core.fp_pipeline.fpiu_unit.queue.valids_3) ||
	  (soc2.core.fp_pipeline.fpiu_unit.queue.value == 3'h4 && soc2.core.fp_pipeline.fpiu_unit.queue.valids_4) ||
	  (soc2.core.fp_pipeline.fpiu_unit.queue.value == 3'h5 && soc2.core.fp_pipeline.fpiu_unit.queue.valids_5) ||
	  (soc2.core.fp_pipeline.fpiu_unit.queue.value == 3'h6 && soc2.core.fp_pipeline.fpiu_unit.queue.valids_6)
	  ?
	  !soc2.core.fp_pipeline.fpiu_unit.queue.do_enq
	  :
	  1'b1
	) &&
	(
	  (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value == 2'h0 && soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0) ||
	  (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value == 2'h1 && soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1) ||
	  (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value == 2'h2 && soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2)
	  ?
	  !soc2.core.fp_pipeline.fpiu_unit.fp_sdq.do_enq
	  :
	  1'b1
	);
	
	wire BranchKillableQueue_pointers_valid_2;
	assign BranchKillableQueue_pointers_valid_2 =
	(soc2.core.jmp_unit.queue.value < 3'h5) && (soc2.core.jmp_unit.queue.value_1 < 3'h5) &&
	(soc2.core.fp_pipeline.fpiu_unit.queue.value < 3'h7) && (soc2.core.fp_pipeline.fpiu_unit.queue.value_1 < 3'h7) &&
	(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value < 2'h3) && (soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 < 2'h3)
	;
	
	wire [5:0] bkq_jmp_rob_idx_2 [4:0];
	assign bkq_jmp_rob_idx_2[0] = soc2.core.jmp_unit.queue.uops_0_rob_idx;
	assign bkq_jmp_rob_idx_2[1] = soc2.core.jmp_unit.queue.uops_1_rob_idx;
	assign bkq_jmp_rob_idx_2[2] = soc2.core.jmp_unit.queue.uops_2_rob_idx;
	assign bkq_jmp_rob_idx_2[3] = soc2.core.jmp_unit.queue.uops_3_rob_idx;
	assign bkq_jmp_rob_idx_2[4] = soc2.core.jmp_unit.queue.uops_4_rob_idx;

	wire bkq_jmp_valids_2 [4:0];
	assign bkq_jmp_valids_2[0] = soc2.core.jmp_unit.queue.valids_0;
	assign bkq_jmp_valids_2[1] = soc2.core.jmp_unit.queue.valids_1;
	assign bkq_jmp_valids_2[2] = soc2.core.jmp_unit.queue.valids_2;
	assign bkq_jmp_valids_2[3] = soc2.core.jmp_unit.queue.valids_3;
	assign bkq_jmp_valids_2[4] = soc2.core.jmp_unit.queue.valids_4;
	  
	wire bkq_jmp_rob_consistency_2;
	assign bkq_jmp_rob_consistency_2 =
	!soc2.core.jmp_unit.queue.io_empty
	?
	  (bkq_jmp_valids_2[(soc2.core.jmp_unit.queue.value_1 + 1) % 5] ? ROBisOlder(bkq_jmp_rob_idx_2[soc2.core.jmp_unit.queue.value_1], bkq_jmp_rob_idx_2[(soc2.core.jmp_unit.queue.value_1 + 1) % 5], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_jmp_valids_2[(soc2.core.jmp_unit.queue.value_1 + 2) % 5] ? ROBisOlder(bkq_jmp_rob_idx_2[(soc2.core.jmp_unit.queue.value_1 + 1) % 5], bkq_jmp_rob_idx_2[(soc2.core.jmp_unit.queue.value_1 + 2) % 5], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_jmp_valids_2[(soc2.core.jmp_unit.queue.value_1 + 3) % 5] ? ROBisOlder(bkq_jmp_rob_idx_2[(soc2.core.jmp_unit.queue.value_1 + 2) % 5], bkq_jmp_rob_idx_2[(soc2.core.jmp_unit.queue.value_1 + 3) % 5], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_jmp_valids_2[(soc2.core.jmp_unit.queue.value_1 + 4) % 5] ? ROBisOlder(bkq_jmp_rob_idx_2[(soc2.core.jmp_unit.queue.value_1 + 3) % 5], bkq_jmp_rob_idx_2[(soc2.core.jmp_unit.queue.value_1 + 4) % 5], soc2.core.rob.io_rob_head_idx) : 1'b1)
	:
	  1'b1;

	wire [5:0] bkq_fp_rob_idx_2 [6:0];
	assign bkq_fp_rob_idx_2[0] = soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx;
	assign bkq_fp_rob_idx_2[1] = soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx;
	assign bkq_fp_rob_idx_2[2] = soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx;
	assign bkq_fp_rob_idx_2[3] = soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx;
	assign bkq_fp_rob_idx_2[4] = soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx;
	assign bkq_fp_rob_idx_2[5] = soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx;
	assign bkq_fp_rob_idx_2[6] = soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx;


	wire bkq_fp_valids_2 [6:0];
	assign bkq_fp_valids_2[0] = soc2.core.fp_pipeline.fpiu_unit.queue.valids_0;
	assign bkq_fp_valids_2[1] = soc2.core.fp_pipeline.fpiu_unit.queue.valids_1;
	assign bkq_fp_valids_2[2] = soc2.core.fp_pipeline.fpiu_unit.queue.valids_2;
	assign bkq_fp_valids_2[3] = soc2.core.fp_pipeline.fpiu_unit.queue.valids_3;
	assign bkq_fp_valids_2[4] = soc2.core.fp_pipeline.fpiu_unit.queue.valids_4;
	assign bkq_fp_valids_2[5] = soc2.core.fp_pipeline.fpiu_unit.queue.valids_5;
	assign bkq_fp_valids_2[6] = soc2.core.fp_pipeline.fpiu_unit.queue.valids_6;

	wire bkq_fp_rob_consistency_2;
	assign bkq_fp_rob_consistency_2 =
	!soc2.core.fp_pipeline.fpiu_unit.queue.io_empty
	?
	  (bkq_fp_valids_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 1) % 7] ? ROBisOlder(bkq_fp_rob_idx_2[soc2.core.fp_pipeline.fpiu_unit.queue.value_1], bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 1) % 7], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 2) % 7] ? ROBisOlder(bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 1) % 7], bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 2) % 7], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 3) % 7] ? ROBisOlder(bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 2) % 7], bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 3) % 7], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 4) % 7] ? ROBisOlder(bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 3) % 7], bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 4) % 7], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 5) % 7] ? ROBisOlder(bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 4) % 7], bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 5) % 7], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_valids_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 6) % 7] ? ROBisOlder(bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 5) % 7], bkq_fp_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.queue.value_1 + 6) % 7], soc2.core.rob.io_rob_head_idx) : 1'b1)
	:
	  1'b1;

	wire [5:0] bkq_fp_1_rob_idx_2 [2:0];
	assign bkq_fp_1_rob_idx_2[0] = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx;
	assign bkq_fp_1_rob_idx_2[1] = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx;
	assign bkq_fp_1_rob_idx_2[2] = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx;

	wire bkq_fp_1_valids_2 [2:0];
	assign bkq_fp_1_valids_2[0] = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0;
	assign bkq_fp_1_valids_2[1] = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1;
	assign bkq_fp_1_valids_2[2] = soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2;
	  
	wire bkq_fp_1_rob_consistency_2;
	assign bkq_fp_1_rob_consistency_2 =
	!soc2.core.fp_pipeline.fpiu_unit.fp_sdq.io_empty
	?
	  (bkq_fp_1_valids_2[(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 1) % 3] ? ROBisOlder(bkq_fp_1_rob_idx_2[soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value_1], bkq_fp_1_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 1) % 3], soc2.core.rob.io_rob_head_idx) : 1'b1) &&
	  (bkq_fp_1_valids_2[(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 2) % 3] ? ROBisOlder(bkq_fp_1_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 1) % 3], bkq_fp_1_rob_idx_2[(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.value_1 + 2) % 3], soc2.core.rob.io_rob_head_idx) : 1'b1)
	:
	  1'b1;

	/*wire ROB_uops_equal_STQ_2;
	assign ROB_uops_equal_STQ_2 =
	  ROB_exists_in_STQ(6'h0, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h1, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h2, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h3, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h4, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h5, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h6, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h7, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h8, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h9, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'ha, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'hb, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'hc, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'hd, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'he, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'hf, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h10, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h11, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h12, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h13, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h14, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h15, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h16, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h17, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h18, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h19, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h1a, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h1b, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h1c, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h1d, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h1e, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h1f, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h20, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h21, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h22, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h23, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h24, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h25, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h26, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h27, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h28, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h29, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h2a, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h2b, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h2c, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h2d, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h2e, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h2f, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h30, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h31, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h32, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h33, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h34, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h35, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h36, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h37, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h38, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h39, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h3a, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h3b, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h3c, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h3d, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h3e, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2) &&
	  ROB_exists_in_STQ(6'h3f, rob_valids_2, rob_uses_stq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, stq_rob_idx_2, rob_stq_indexes_2, stq_valids_2, stq_committed_2);

	wire ROB_uops_equal_LDQ_2;
	assign ROB_uops_equal_LDQ_2 =
	  ROB_exists_in_LDQ(6'h0, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h1, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h2, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h3, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h4, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h5, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h6, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h7, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h8, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h9, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'ha, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'hb, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'hc, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'hd, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'he, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'hf, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h10, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h11, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h12, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h13, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h14, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h15, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h16, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h17, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h18, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h19, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h1a, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h1b, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h1c, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h1d, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h1e, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h1f, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h20, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h21, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h22, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h23, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h24, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h25, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h26, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h27, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h28, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h29, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h2a, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h2b, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h2c, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h2d, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h2e, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h2f, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h30, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h31, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h32, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h33, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h34, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h35, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h36, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h37, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h38, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h39, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h3a, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h3b, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h3c, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h3d, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h3e, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2) &&
	  ROB_exists_in_LDQ(6'h3f, rob_valids_2, rob_uses_ldq_2, soc2.core.rob.rob_state, soc2.core.rob.REG_1, rob_exception_2, ldq_rob_idx_2, rob_ldq_indexes_2, ldq_valids_2);*/

	wire STQ_uops_equals_ROB_2;
	assign STQ_uops_equals_ROB_2 =
	  STQ_exists_in_ROB(4'h0, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'h1, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'h2, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'h3, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'h4, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'h5, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'h6, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'h7, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'h8, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'h9, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'ha, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'hb, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'hc, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'hd, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'he, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2) &&
	  STQ_exists_in_ROB(4'hf, stq_valids_2, stq_committed_2, rob_uses_stq_2, stq_rob_idx_2, rob_valids_2);

	wire LDQ_uops_equals_ROB_2;
	assign LDQ_uops_equals_ROB_2 =
	  LDQ_exists_in_ROB(4'h0, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'h1, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'h2, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'h3, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'h4, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'h5, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'h6, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'h7, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'h8, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'h9, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'ha, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'hb, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'hc, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'hd, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'he, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2) &&
	  LDQ_exists_in_ROB(4'hf, ldq_valids_2, rob_uses_ldq_2, ldq_rob_idx_2, rob_valids_2);


	wire ldq_uses_ldq_2[15:0];
	assign ldq_uses_ldq_2[0] = soc2.lsu.ldq_0_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[1] = soc2.lsu.ldq_1_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[2] = soc2.lsu.ldq_2_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[3] = soc2.lsu.ldq_3_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[4] = soc2.lsu.ldq_4_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[5] = soc2.lsu.ldq_5_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[6] = soc2.lsu.ldq_6_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[7] = soc2.lsu.ldq_7_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[8] = soc2.lsu.ldq_8_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[9] = soc2.lsu.ldq_9_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[10] = soc2.lsu.ldq_10_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[11] = soc2.lsu.ldq_11_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[12] = soc2.lsu.ldq_12_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[13] = soc2.lsu.ldq_13_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[14] = soc2.lsu.ldq_14_bits_uop_uses_ldq;
	assign ldq_uses_ldq_2[15] = soc2.lsu.ldq_15_bits_uop_uses_ldq;

	wire stq_uses_stq_2[15:0];
	assign stq_uses_stq_2[0] = soc2.lsu.stq_0_bits_uop_uses_stq;
	assign stq_uses_stq_2[1] = soc2.lsu.stq_1_bits_uop_uses_stq;
	assign stq_uses_stq_2[2] = soc2.lsu.stq_2_bits_uop_uses_stq;
	assign stq_uses_stq_2[3] = soc2.lsu.stq_3_bits_uop_uses_stq;
	assign stq_uses_stq_2[4] = soc2.lsu.stq_4_bits_uop_uses_stq;
	assign stq_uses_stq_2[5] = soc2.lsu.stq_5_bits_uop_uses_stq;
	assign stq_uses_stq_2[6] = soc2.lsu.stq_6_bits_uop_uses_stq;
	assign stq_uses_stq_2[7] = soc2.lsu.stq_7_bits_uop_uses_stq;
	assign stq_uses_stq_2[8] = soc2.lsu.stq_8_bits_uop_uses_stq;
	assign stq_uses_stq_2[9] = soc2.lsu.stq_9_bits_uop_uses_stq;
	assign stq_uses_stq_2[10] = soc2.lsu.stq_10_bits_uop_uses_stq;
	assign stq_uses_stq_2[11] = soc2.lsu.stq_11_bits_uop_uses_stq;
	assign stq_uses_stq_2[12] = soc2.lsu.stq_12_bits_uop_uses_stq;
	assign stq_uses_stq_2[13] = soc2.lsu.stq_13_bits_uop_uses_stq;
	assign stq_uses_stq_2[14] = soc2.lsu.stq_14_bits_uop_uses_stq;
	assign stq_uses_stq_2[15] = soc2.lsu.stq_15_bits_uop_uses_stq;

	wire buffers_equal_ROB_2;
	assign buffers_equal_ROB_2 =
	Buffer_exists_in_ROB_stq_idx_only(soc2.core.b2_mispredict, stq_committed_2, soc2.core.b2_uop_stq_idx, rob_valids_2, soc2.core.b2_uop_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc2.core.brinfos_0_valid, stq_committed_2, soc2.core.brinfos_0_uop_stq_idx, rob_valids_2, soc2.core.brinfos_0_uop_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc2.core.brinfos_1_valid, stq_committed_2, soc2.core.brinfos_1_uop_stq_idx, rob_valids_2, soc2.core.brinfos_1_uop_rob_idx) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.csr_exe_unit.alu.r_valids_0, soc2.core.csr_exe_unit.alu.r_uops_0_uses_stq, rob_valids_2, soc2.core.csr_exe_unit.alu.r_uops_0_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq((soc2.core.csr_exe_unit.div.div.state == 3'h3) || (soc2.core.csr_exe_unit.div.div.state == 3'h7), soc2.core.csr_exe_unit.div.r_uop_uses_stq, rob_valids_2, soc2.core.csr_exe_unit.div.r_uop_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_0.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_0.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_1.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_1.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_2.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_2.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_3.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_3.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_4.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_4.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_5.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_5.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_6.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_6.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_7.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_7.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_8.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_8.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_9.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_9.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_10.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_10.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_11.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_11.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_12.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_12.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_13.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_13.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_14.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_14.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fp_issue_unit.slots_15.io_valid, soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fp_issue_unit.slots_15.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.queue.valids_0, soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_0_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.queue.valids_1, soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_1_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.queue.valids_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_2_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.queue.valids_3, soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_3_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.queue.valids_4, soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_4_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.queue.valids_5, soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_5_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.queue.valids_6, soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.queue.uops_6_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_0, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_0_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_1, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_1_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.fp_pipeline.fpiu_unit.fp_sdq.valids_2, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fp_sdq.uops_2_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_no_idx(soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_val, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_uses_stq, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_buffer_req_uop_uses_ldq) &&
	Buffer_exists_in_ROB_no_idx(soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_uses_stq, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_uop_uses_ldq) &&
	Buffer_exists_in_ROB_no_idx(soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_val, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_uses_stq, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_out_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_0, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_0_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_1, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_1_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_2_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fpiu_unit.fpu.r_valids_3, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.fp_pipeline.fpiu_unit.fpu.r_uops_3_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fregister_read.exe_reg_valids_0, soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_rob_idx, rob_uses_stq_2, rob_uses_ldq_2,soc2.core.fp_pipeline.fregister_read.exe_reg_uops_0_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.fp_pipeline.fregister_read.rrd_valids_0_REG, soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uses_stq, stq_committed_2, soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_stq_idx, rob_valids_2, soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_rob_idx, rob_uses_stq_2, rob_uses_ldq_2,soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_0.io_valid, soc2.core.int_issue_unit.slots_0.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_0.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_0.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_0.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_1.io_valid, soc2.core.int_issue_unit.slots_1.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_1.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_1.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_1.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_2.io_valid, soc2.core.int_issue_unit.slots_2.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_2.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_2.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_2.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_3.io_valid, soc2.core.int_issue_unit.slots_3.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_3.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_3.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_3.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_4.io_valid, soc2.core.int_issue_unit.slots_4.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_4.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_4.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_4.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_5.io_valid, soc2.core.int_issue_unit.slots_5.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_5.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_5.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_5.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_6.io_valid, soc2.core.int_issue_unit.slots_6.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_6.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_6.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_6.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_7.io_valid, soc2.core.int_issue_unit.slots_7.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_7.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_7.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_7.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_8.io_valid, soc2.core.int_issue_unit.slots_8.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_8.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_8.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_8.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_9.io_valid, soc2.core.int_issue_unit.slots_9.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_9.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_9.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_9.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_10.io_valid, soc2.core.int_issue_unit.slots_10.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_10.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_10.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_10.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_11.io_valid, soc2.core.int_issue_unit.slots_11.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_11.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_11.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_11.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_12.io_valid, soc2.core.int_issue_unit.slots_12.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_12.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_12.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_12.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_13.io_valid, soc2.core.int_issue_unit.slots_13.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_13.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_13.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_13.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_14.io_valid, soc2.core.int_issue_unit.slots_14.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_14.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_14.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_14.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_15.io_valid, soc2.core.int_issue_unit.slots_15.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_15.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_15.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_15.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_16.io_valid, soc2.core.int_issue_unit.slots_16.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_16.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_16.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_16.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_17.io_valid, soc2.core.int_issue_unit.slots_17.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_17.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_17.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_17.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_18.io_valid, soc2.core.int_issue_unit.slots_18.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_18.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_18.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_18.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.int_issue_unit.slots_19.io_valid, soc2.core.int_issue_unit.slots_19.slot_uop_uses_stq, stq_committed_2, soc2.core.int_issue_unit.slots_19.slot_uop_stq_idx, rob_valids_2, soc2.core.int_issue_unit.slots_19.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.int_issue_unit.slots_19.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.iregister_read.exe_reg_valids_0, soc2.core.iregister_read.exe_reg_uops_0_uses_stq, stq_committed_2, soc2.core.iregister_read.exe_reg_uops_0_stq_idx, rob_valids_2, soc2.core.iregister_read.exe_reg_uops_0_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.iregister_read.exe_reg_uops_0_uses_ldq) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.iregister_read.exe_reg_valids_1, soc2.core.iregister_read.exe_reg_uops_1_uses_stq, stq_committed_2, soc2.core.iregister_read.exe_reg_uops_1_stq_idx, rob_valids_2, soc2.core.iregister_read.exe_reg_uops_1_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.iregister_read.exe_reg_valids_2, soc2.core.iregister_read.exe_reg_uops_2_uses_stq, stq_committed_2, soc2.core.iregister_read.exe_reg_uops_2_stq_idx, rob_valids_2, soc2.core.iregister_read.exe_reg_uops_2_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB(soc2.core.iregister_read.rrd_valids_0_REG, soc2.core.iregister_read.rrd_uops_0_REG_uses_stq, stq_committed_2, soc2.core.iregister_read.rrd_uops_0_REG_stq_idx, rob_valids_2, soc2.core.iregister_read.rrd_uops_0_REG_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.iregister_read.rrd_uops_0_REG_uses_ldq) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.iregister_read.rrd_valids_1_REG, soc2.core.iregister_read.rrd_uops_1_REG_uses_stq, stq_committed_2, soc2.core.iregister_read.rrd_uops_1_REG_stq_idx, rob_valids_2, soc2.core.iregister_read.rrd_uops_1_REG_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_stq(soc2.core.iregister_read.rrd_valids_2_REG, soc2.core.iregister_read.rrd_uops_2_REG_uses_stq, stq_committed_2, soc2.core.iregister_read.rrd_uops_2_REG_stq_idx, rob_valids_2, soc2.core.iregister_read.rrd_uops_2_REG_rob_idx, rob_uses_stq_2) &&
	//(soc2.core.jmp_unit.queue.ram_fflags_valid ? rob_valids_2[soc2.core.jmp_unit.queue.ram_fflags_bits_uop_rob_idx] : 1'b1) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.queue.valids_0, soc2.core.jmp_unit.queue.uops_0_uses_stq, rob_valids_2, soc2.core.jmp_unit.queue.uops_0_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.queue.valids_1, soc2.core.jmp_unit.queue.uops_1_uses_stq, rob_valids_2, soc2.core.jmp_unit.queue.uops_1_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.queue.valids_2, soc2.core.jmp_unit.queue.uops_2_uses_stq, rob_valids_2, soc2.core.jmp_unit.queue.uops_2_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.queue.valids_3, soc2.core.jmp_unit.queue.uops_3_uses_stq, rob_valids_2, soc2.core.jmp_unit.queue.uops_3_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.queue.valids_4, soc2.core.jmp_unit.queue.uops_4_uses_stq, rob_valids_2, soc2.core.jmp_unit.queue.uops_4_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.alu.r_valids_0, soc2.core.jmp_unit.alu.r_uops_0_uses_stq, rob_valids_2, soc2.core.jmp_unit.alu.r_uops_0_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.alu.r_valids_1, soc2.core.jmp_unit.alu.r_uops_1_uses_stq, rob_valids_2, soc2.core.jmp_unit.alu.r_uops_1_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.alu.r_valids_2, soc2.core.jmp_unit.alu.r_uops_2_uses_stq, rob_valids_2, soc2.core.jmp_unit.alu.r_uops_2_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.ifpu.r_valids_0, soc2.core.jmp_unit.ifpu.r_uops_0_uses_stq, rob_valids_2, soc2.core.jmp_unit.ifpu.r_uops_0_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.ifpu.r_valids_1, soc2.core.jmp_unit.ifpu.r_uops_1_uses_stq, rob_valids_2, soc2.core.jmp_unit.ifpu.r_uops_1_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.imul.r_valids_0, soc2.core.jmp_unit.imul.r_uops_0_uses_stq, rob_valids_2, soc2.core.jmp_unit.imul.r_uops_0_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.imul.r_valids_1, soc2.core.jmp_unit.imul.r_uops_1_uses_stq, rob_valids_2, soc2.core.jmp_unit.imul.r_uops_1_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB_only_uses_stq(soc2.core.jmp_unit.imul.r_valids_2, soc2.core.jmp_unit.imul.r_uops_2_uses_stq, rob_valids_2, soc2.core.jmp_unit.imul.r_uops_2_rob_idx, rob_uses_stq_2) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_0.io_valid, soc2.core.mem_issue_unit.slots_0.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_0.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_0.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_0.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_1.io_valid, soc2.core.mem_issue_unit.slots_1.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_1.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_1.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_1.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_2.io_valid, soc2.core.mem_issue_unit.slots_2.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_2.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_2.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_2.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_3.io_valid, soc2.core.mem_issue_unit.slots_3.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_3.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_3.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_3.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_4.io_valid, soc2.core.mem_issue_unit.slots_4.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_4.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_4.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_4.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_5.io_valid, soc2.core.mem_issue_unit.slots_5.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_5.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_5.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_5.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_6.io_valid, soc2.core.mem_issue_unit.slots_6.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_6.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_6.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_6.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_7.io_valid, soc2.core.mem_issue_unit.slots_7.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_7.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_7.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_7.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_8.io_valid, soc2.core.mem_issue_unit.slots_8.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_8.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_8.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_8.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_9.io_valid, soc2.core.mem_issue_unit.slots_9.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_9.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_9.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_9.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_10.io_valid, soc2.core.mem_issue_unit.slots_10.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_10.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_10.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_10.slot_uop_uses_ldq) &&
	Buffer_exists_in_ROB(soc2.core.mem_issue_unit.slots_11.io_valid, soc2.core.mem_issue_unit.slots_11.slot_uop_uses_stq, stq_committed_2, soc2.core.mem_issue_unit.slots_11.slot_uop_stq_idx, rob_valids_2, soc2.core.mem_issue_unit.slots_11.slot_uop_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.core.mem_issue_unit.slots_11.slot_uop_uses_ldq) &&
	(soc2.core.rob.r_xcpt_val ? rob_valids_2[soc2.core.rob.r_xcpt_uop_rob_idx] : 1'b1) &&
	//Buffer_exists_in_LDQ(soc2.dcache.s1_valid_0, soc2.dcache.s1_req_0_uop_uses_ldq, ldq_valids_2, soc2.dcache.s1_req_0_uop_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.s1_valid_0 && (soc2.dcache.s1_type != 3'b0 || soc2.dcache.s1_req_0_uop_is_amo), soc2.dcache.s1_req_0_uop_uses_stq, stq_valids_2, soc2.dcache.s1_req_0_uop_stq_idx, stq_uses_stq_2) &&
	//Buffer_exists_in_LDQ(soc2.dcache.s2_valid_0, soc2.dcache.s2_req_0_uop_uses_ldq, ldq_valids_2, soc2.dcache.s2_req_0_uop_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.s2_valid_0 && (soc2.dcache.s2_type != 3'b0 || soc2.dcache.s2_req_0_uop_is_amo), soc2.dcache.s2_req_0_uop_uses_stq, stq_valids_2, soc2.dcache.s2_req_0_uop_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mmios_0.state != 2'b0, soc2.dcache.mshrs.mmios_0.req_uop_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mmios_0.req_uop_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(!soc2.dcache.mshrs.mmios_0.io_req_valid, soc2.dcache.mshrs.mmios_0.req_uop_uses_stq, stq_valids_2, soc2.dcache.mshrs.mmios_0.req_uop_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_0, soc2.dcache.mshrs.mshrs_0.rpq.uops_0_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_0_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_0, soc2.dcache.mshrs.mshrs_0.rpq.uops_0_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_0_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_1, soc2.dcache.mshrs.mshrs_0.rpq.uops_1_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_1_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_1, soc2.dcache.mshrs.mshrs_0.rpq.uops_1_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_1_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_2_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_2_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_2_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_2_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_3, soc2.dcache.mshrs.mshrs_0.rpq.uops_3_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_3_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_3, soc2.dcache.mshrs.mshrs_0.rpq.uops_3_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_3_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_4, soc2.dcache.mshrs.mshrs_0.rpq.uops_4_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_4_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_4, soc2.dcache.mshrs.mshrs_0.rpq.uops_4_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_4_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_5, soc2.dcache.mshrs.mshrs_0.rpq.uops_5_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_5_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_5, soc2.dcache.mshrs.mshrs_0.rpq.uops_5_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_5_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_6, soc2.dcache.mshrs.mshrs_0.rpq.uops_6_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_6_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_6, soc2.dcache.mshrs.mshrs_0.rpq.uops_6_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_6_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_7, soc2.dcache.mshrs.mshrs_0.rpq.uops_7_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_7_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_7, soc2.dcache.mshrs.mshrs_0.rpq.uops_7_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_7_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_8, soc2.dcache.mshrs.mshrs_0.rpq.uops_8_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_8_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_8, soc2.dcache.mshrs.mshrs_0.rpq.uops_8_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_8_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_9, soc2.dcache.mshrs.mshrs_0.rpq.uops_9_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_9_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_9, soc2.dcache.mshrs.mshrs_0.rpq.uops_9_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_9_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_10, soc2.dcache.mshrs.mshrs_0.rpq.uops_10_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_10_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_10, soc2.dcache.mshrs.mshrs_0.rpq.uops_10_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_10_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_11, soc2.dcache.mshrs.mshrs_0.rpq.uops_11_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_11_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_11, soc2.dcache.mshrs.mshrs_0.rpq.uops_11_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_11_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_12, soc2.dcache.mshrs.mshrs_0.rpq.uops_12_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_12_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_12, soc2.dcache.mshrs.mshrs_0.rpq.uops_12_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_12_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_13, soc2.dcache.mshrs.mshrs_0.rpq.uops_13_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_13_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_13, soc2.dcache.mshrs.mshrs_0.rpq.uops_13_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_13_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_14, soc2.dcache.mshrs.mshrs_0.rpq.uops_14_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_14_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_14, soc2.dcache.mshrs.mshrs_0.rpq.uops_14_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_14_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_15, soc2.dcache.mshrs.mshrs_0.rpq.uops_15_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_15_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_0.rpq.valids_15, soc2.dcache.mshrs.mshrs_0.rpq.uops_15_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_0.rpq.uops_15_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_0, soc2.dcache.mshrs.mshrs_1.rpq.uops_0_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_0_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_0, soc2.dcache.mshrs.mshrs_1.rpq.uops_0_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_0_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_1, soc2.dcache.mshrs.mshrs_1.rpq.uops_1_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_1_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_1, soc2.dcache.mshrs.mshrs_1.rpq.uops_1_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_1_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_2_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_2_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_2_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_2_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_3, soc2.dcache.mshrs.mshrs_1.rpq.uops_3_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_3_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_3, soc2.dcache.mshrs.mshrs_1.rpq.uops_3_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_3_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_4, soc2.dcache.mshrs.mshrs_1.rpq.uops_4_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_4_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_4, soc2.dcache.mshrs.mshrs_1.rpq.uops_4_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_4_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_5, soc2.dcache.mshrs.mshrs_1.rpq.uops_5_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_5_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_5, soc2.dcache.mshrs.mshrs_1.rpq.uops_5_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_5_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_6, soc2.dcache.mshrs.mshrs_1.rpq.uops_6_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_6_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_6, soc2.dcache.mshrs.mshrs_1.rpq.uops_6_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_6_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_7, soc2.dcache.mshrs.mshrs_1.rpq.uops_7_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_7_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_7, soc2.dcache.mshrs.mshrs_1.rpq.uops_7_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_7_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_8, soc2.dcache.mshrs.mshrs_1.rpq.uops_8_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_8_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_8, soc2.dcache.mshrs.mshrs_1.rpq.uops_8_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_8_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_9, soc2.dcache.mshrs.mshrs_1.rpq.uops_9_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_9_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_9, soc2.dcache.mshrs.mshrs_1.rpq.uops_9_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_9_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_10, soc2.dcache.mshrs.mshrs_1.rpq.uops_10_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_10_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_10, soc2.dcache.mshrs.mshrs_1.rpq.uops_10_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_10_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_11, soc2.dcache.mshrs.mshrs_1.rpq.uops_11_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_11_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_11, soc2.dcache.mshrs.mshrs_1.rpq.uops_11_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_11_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_12, soc2.dcache.mshrs.mshrs_1.rpq.uops_12_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_12_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_12, soc2.dcache.mshrs.mshrs_1.rpq.uops_12_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_12_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_13, soc2.dcache.mshrs.mshrs_1.rpq.uops_13_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_13_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_13, soc2.dcache.mshrs.mshrs_1.rpq.uops_13_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_13_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_14, soc2.dcache.mshrs.mshrs_1.rpq.uops_14_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_14_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_14, soc2.dcache.mshrs.mshrs_1.rpq.uops_14_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_14_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_15, soc2.dcache.mshrs.mshrs_1.rpq.uops_15_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_15_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.mshrs_1.rpq.valids_15, soc2.dcache.mshrs.mshrs_1.rpq.uops_15_uses_stq, stq_valids_2, soc2.dcache.mshrs.mshrs_1.rpq.uops_15_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.respq.valids_0, soc2.dcache.mshrs.respq.uops_0_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.respq.uops_0_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.respq.valids_0, soc2.dcache.mshrs.respq.uops_0_uses_stq, stq_valids_2, soc2.dcache.mshrs.respq.uops_0_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.respq.valids_1, soc2.dcache.mshrs.respq.uops_1_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.respq.uops_1_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.respq.valids_1, soc2.dcache.mshrs.respq.uops_1_uses_stq, stq_valids_2, soc2.dcache.mshrs.respq.uops_1_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.respq.valids_2, soc2.dcache.mshrs.respq.uops_2_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.respq.uops_2_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.respq.valids_2, soc2.dcache.mshrs.respq.uops_2_uses_stq, stq_valids_2, soc2.dcache.mshrs.respq.uops_2_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_LDQ(soc2.dcache.mshrs.respq.valids_3, soc2.dcache.mshrs.respq.uops_3_uses_ldq, ldq_valids_2, soc2.dcache.mshrs.respq.uops_3_ldq_idx, ldq_uses_ldq_2) &&
	//Buffer_exists_in_STQ(soc2.dcache.mshrs.respq.valids_3, soc2.dcache.mshrs.respq.uops_3_uses_stq, stq_valids_2, soc2.dcache.mshrs.respq.uops_3_stq_idx, stq_uses_stq_2) &&
	Buffer_exists_in_ROB_stq_idx_only(soc2.lsu.fired_sfence_0 || soc2.lsu.fired_load_incoming_REG || soc2.lsu.fired_sta_incoming_REG || soc2.lsu.fired_stad_incoming_REG || soc2.lsu.fired_std_incoming_REG, stq_committed_2, soc2.lsu.mem_incoming_uop_0_stq_idx, rob_valids_2, soc2.lsu.mem_incoming_uop_0_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc2.lsu.fired_stdf_incoming, stq_committed_2, soc2.lsu.mem_stdf_uop_stq_idx, rob_valids_2, soc2.lsu.mem_stdf_uop_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc2.lsu.fired_sta_incoming_REG || soc2.lsu.fired_stad_incoming_REG || soc2.lsu.fired_std_incoming_REG, stq_committed_2, soc2.lsu.mem_stq_incoming_e_0_bits_uop_stq_idx, rob_valids_2, soc2.lsu.mem_stq_incoming_e_0_bits_uop_rob_idx) &&
	Buffer_exists_in_ROB_stq_idx_only(soc2.lsu.fired_sta_retry_REG, stq_committed_2, soc2.lsu.mem_stq_retry_e_bits_uop_stq_idx, rob_valids_2, soc2.lsu.mem_stq_retry_e_bits_uop_rob_idx) &&
	Buffer_exists_in_ROB(soc2.lsu.mem_xcpt_valids_0, soc2.lsu.mem_xcpt_uops_0_uses_stq, stq_committed_2, soc2.lsu.mem_xcpt_uops_0_stq_idx, rob_valids_2, soc2.lsu.mem_xcpt_uops_0_rob_idx, rob_uses_stq_2, rob_uses_ldq_2, soc2.lsu.mem_xcpt_uops_0_uses_ldq)
	;
	
	/*
	wire unique_stq_idx_2;
	assign unique_stq_idx_2 = check_uniqueness_stq_idx(rob_valids_2, rob_uses_stq_2, rob_stq_indexes_2);*/
	
	wire stdf_clr_bsy_uses_stq_2;
	assign stdf_clr_bsy_uses_stq_2 = soc2.lsu.stdf_clr_bsy_valid ? rob_uses_stq_2[soc2.lsu.stdf_clr_bsy_rob_idx] : 1'b1;

	wire fdivsqrt_consistency_2;
	assign fdivsqrt_consistency_2 =
	(soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.r_divsqrt_val
	?
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A != 3'b0
	  ?
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B == 4'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C == 3'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E == 3'b0)
	  :
	    1'b1
	  ) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B != 4'b0
	  ?
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A == 3'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C == 3'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E == 3'b0)
	  :
	    1'b1
	  ) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C != 3'b0
	  ?
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B == 4'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A == 3'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E == 3'b0)
	  :
	    1'b1
	  ) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E != 3'b0
	  ?
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B == 4'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C == 3'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A == 3'b0)
	  :
	    1'b1
	  ) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PA
	  ?
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PB == 1'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PC == 1'b0)
	  :
	    1'b1
	  ) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PB
	  ?
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PA == 1'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PC == 1'b0)
	  :
	    1'b1
	  ) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PC
	  ?
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PB == 1'b0) &&
	    (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PA == 1'b0)
	  :
	    1'b1
	  )
	:
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_A == 3'b0) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_B == 4'b0) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_C == 3'b0) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.cycleNum_E == 3'b0) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PA == 1'b0) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PB == 1'b0) &&
	  (soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.divsqrt.ds.divSqrtRecF64ToRaw.valid_PC == 1'b0)
	);
	
	wire unique_write_port_addr_2;
	assign unique_write_port_addr_2 =
		(soc2.core.iregfile.io_write_ports_0_valid && soc2.core.iregfile.io_write_ports_1_valid ? soc2.core.iregfile.io_write_ports_0_bits_addr != soc2.core.iregfile.io_write_ports_1_bits_addr : 1'b1) &&
		(soc2.core.iregfile.io_write_ports_0_valid && soc2.core.iregfile.io_write_ports_2_valid ? soc2.core.iregfile.io_write_ports_0_bits_addr != soc2.core.iregfile.io_write_ports_2_bits_addr : 1'b1) &&
		(soc2.core.iregfile.io_write_ports_1_valid && soc2.core.iregfile.io_write_ports_2_valid ? soc2.core.iregfile.io_write_ports_1_bits_addr != soc2.core.iregfile.io_write_ports_2_bits_addr : 1'b1)
	;
	
	wire lsu_req_consistent_2;
	assign lsu_req_consistent_2 =
		soc2.lsu.io_core_exe_0_req_valid
		?
			(soc2.lsu.io_core_exe_0_req_bits_uop_ctrl_is_load == soc2.lsu.io_core_exe_0_req_bits_uop_uses_ldq) &&
			((soc2.lsu.io_core_exe_0_req_bits_uop_ctrl_is_sta || soc2.lsu.io_core_exe_0_req_bits_uop_ctrl_is_std) == soc2.lsu.io_core_exe_0_req_bits_uop_uses_stq)
		:
			1'b1;
			
	wire csr_req_not_speculative_2;
	assign csr_req_not_speculative_2 = soc2.core.csr_exe_unit.io_req_valid && soc2.core.csr_exe_unit.io_req_bits_uop_ctrl_csr_cmd != 3'b0 ? soc2.core.csr_exe_unit.io_req_bits_uop_br_mask == 12'b0 : 1'b1;
	
	wire lsu_req_uses_queue_2;
	assign lsu_req_uses_queue_2 = soc2.lsu.io_core_exe_0_req_valid ? soc2.lsu.io_core_exe_0_req_bits_uop_uses_ldq || soc2.lsu.io_core_exe_0_req_bits_uop_uses_stq || (soc2.lsu.io_core_exe_0_req_bits_sfence_valid && soc2.lsu.io_core_exe_0_req_bits_uop_br_mask == 12'b0): 1'b1;
	
	wire dmem_resp_amo_2;
	assign dmem_resp_amo_2 =
	soc2.lsu.io_dmem_resp_0_valid && soc2.lsu.io_dmem_resp_0_bits_uop_is_amo
	?
		soc2.lsu.io_dmem_resp_0_bits_uop_uses_stq && stq_valids_2[soc2.lsu.io_dmem_resp_0_bits_uop_stq_idx] &&
		(rob_branch_masks_2[stq_rob_idx_2[soc2.lsu.io_dmem_resp_0_bits_uop_stq_idx]] == 12'b0) &&
		!stq_committed_2[soc2.lsu.io_dmem_resp_0_bits_uop_stq_idx] &&
		soc2.lsu.stq_head == soc2.lsu.io_dmem_resp_0_bits_uop_stq_idx &&
		soc2.core.rob.io_rob_head_idx == stq_rob_idx_2[soc2.lsu.io_dmem_resp_0_bits_uop_stq_idx] &&
		soc2.core.rob.io_rob_tail_idx == ((stq_rob_idx_2[soc2.lsu.io_dmem_resp_0_bits_uop_stq_idx] + 1) % 64)
	:
		1'b1
	;
	
	wire buffers_equal_STQ_2;
	assign buffers_equal_STQ_2 = 
		(soc2.lsu.fired_stdf_incoming && !stq_committed_2[soc2.lsu.mem_stdf_uop_stq_idx] ? stq_valids_2[soc2.lsu.mem_stdf_uop_stq_idx] && soc2.lsu.mem_stdf_uop_rob_idx == stq_rob_idx_2[soc2.lsu.mem_stdf_uop_stq_idx] : 1'b1) &&
		(soc2.core.iregister_read.exe_reg_valids_0 && soc2.core.iregister_read.exe_reg_uops_0_uses_stq && !stq_committed_2[soc2.core.iregister_read.exe_reg_uops_0_stq_idx] ? stq_valids_2[soc2.core.iregister_read.exe_reg_uops_0_stq_idx] && soc2.core.iregister_read.exe_reg_uops_0_rob_idx == stq_rob_idx_2[soc2.core.iregister_read.exe_reg_uops_0_stq_idx] : 1'b1);
	
	wire buffers_equal_LDQ_2;
	assign buffers_equal_LDQ_2 =
	  (soc2.core.iregister_read.exe_reg_valids_0 && soc2.core.iregister_read.exe_reg_uops_0_uses_ldq ? ldq_valids_2[soc2.core.iregister_read.exe_reg_uops_0_ldq_idx] && soc2.core.iregister_read.exe_reg_uops_0_rob_idx == ldq_rob_idx_2[soc2.core.iregister_read.exe_reg_uops_0_ldq_idx] : 1'b1);

	
	wire ldq_head_empty_2;
	assign ldq_head_empty_2 = !ldq_valids_2[soc2.lsu.ldq_head] == (!ldq_valids_2[0] && !ldq_valids_2[1] && !ldq_valids_2[2] && !ldq_valids_2[3] && !ldq_valids_2[4] && !ldq_valids_2[5] && !ldq_valids_2[6] && !ldq_valids_2[7] && !ldq_valids_2[8] &&
	 !ldq_valids_2[9] && !ldq_valids_2[10] && !ldq_valids_2[11] && !ldq_valids_2[12] && !ldq_valids_2[13] && !ldq_valids_2[14] && !ldq_valids_2[15]);

	wire unique_ldq_rob_idx_2;
	assign unique_ldq_rob_idx_2 = check_uniqueness_ldq_rob_idx(ldq_valids_2, ldq_rob_idx_2);	
	
	/*wire mem_xcpt_consistency_2;
	assign mem_xcpt_consistency_2 =
	  soc2.lsu.will_fire_store_commit_0 && soc2.lsu.mem_xcpt_valids_0
	  ?
	    soc2.lsu.mem_xcpt_uops_0_stq_idx == soc2.lsu.stq_execute_head && soc2.lsu.mem_xcpt_uops_0_uses_stq
	  :
	    1'b1;*/
	    
	wire fired_load_incoming_conflicts_2;
	assign fired_load_incoming_conflicts_2 =
	  !(soc2.lsu.fired_load_incoming_REG && soc2.lsu.fired_stad_incoming_REG) &&
	  !(soc2.lsu.fired_load_incoming_REG && soc2.lsu.fired_sta_incoming_REG) &&
	  !(soc2.lsu.fired_load_incoming_REG && soc2.lsu.fired_sfence_0) &&
	  !(soc2.lsu.fired_load_incoming_REG && soc2.lsu.fired_load_retry_REG) &&
	  !(soc2.lsu.fired_load_incoming_REG && soc2.lsu.fired_sta_retry_REG) &&
	  !(soc2.lsu.fired_load_incoming_REG && soc2.lsu.fired_release_0) &&
	  !(soc2.lsu.fired_load_incoming_REG && soc2.lsu.fired_load_wakeup_REG);
	  
	wire fired_stad_incoming_conflicts_2;
	assign fired_stad_incoming_conflicts_2 =
	  !(soc2.lsu.fired_stad_incoming_REG && soc2.lsu.fired_sta_incoming_REG) &&
	  !(soc2.lsu.fired_stad_incoming_REG && soc2.lsu.fired_std_incoming_REG) &&
	  !(soc2.lsu.fired_stad_incoming_REG && soc2.lsu.fired_sfence_0) &&
	  !(soc2.lsu.fired_stad_incoming_REG && soc2.lsu.fired_release_0) &&
	  !(soc2.lsu.fired_stad_incoming_REG && soc2.lsu.fired_load_retry_REG) &&
	  !(soc2.lsu.fired_stad_incoming_REG && soc2.lsu.fired_sta_retry_REG) &&
	  !(soc2.lsu.fired_stad_incoming_REG && soc2.lsu.fired_load_wakeup_REG);

	wire fired_sta_incoming_conflicts_2;
	assign fired_sta_incoming_conflicts_2 =
	  !(soc2.lsu.fired_sta_incoming_REG && soc2.lsu.fired_std_incoming_REG) &&
	  !(soc2.lsu.fired_sta_incoming_REG && soc2.lsu.fired_sfence_0) &&
	  !(soc2.lsu.fired_sta_incoming_REG && soc2.lsu.fired_release_0) &&
	  !(soc2.lsu.fired_sta_incoming_REG && soc2.lsu.fired_load_retry_REG) &&
	  !(soc2.lsu.fired_sta_incoming_REG && soc2.lsu.fired_sta_retry_REG) &&
	  !(soc2.lsu.fired_sta_incoming_REG && soc2.lsu.fired_load_wakeup_REG);

	wire fired_std_incoming_conflicts_2;
	assign fired_std_incoming_conflicts_2 =
	  !(soc2.lsu.fired_std_incoming_REG && soc2.lsu.fired_sfence_0) &&
	  !(soc2.lsu.fired_std_incoming_REG && soc2.lsu.fired_sta_retry_REG);

	wire fired_std_conflicts_2;
	assign fired_std_conflicts_2 = 1'b1;

	wire fired_sfence_conflicts_2;
	assign fired_sfence_conflicts_2 = 
	  !(soc2.lsu.fired_sfence_0 && soc2.lsu.fired_load_retry_REG) &&
	  !(soc2.lsu.fired_sfence_0 && soc2.lsu.fired_sta_retry_REG);

	wire fired_release_conflicts_2;
	assign fired_release_conflicts_2 = 
	  !(soc2.lsu.fired_release_0 && soc2.lsu.fired_load_retry_REG) &&
	  !(soc2.lsu.fired_release_0 && soc2.lsu.fired_sta_retry_REG);

	wire fired_load_retry_conflicts_2;
	assign fired_load_retry_conflicts_2 = 
	  !(soc2.lsu.fired_load_retry_REG && soc2.lsu.fired_sta_retry_REG) &&
	  !(soc2.lsu.fired_load_retry_REG && soc2.lsu.fired_load_wakeup_REG);

	wire fired_sta_retry_conflicts_2;
	assign fired_sta_retry_conflicts_2 = 
	  !(soc2.lsu.fired_sta_retry_REG && soc2.lsu.fired_load_wakeup_REG);
	  
	wire rrd_lrs_types_2;
	assign rrd_lrs_types_2 =
	check_uopc_lrs1_lrs2(soc2.core.iregister_read.rrd_uops_0_REG_uopc, soc2.core.iregister_read.rrd_uops_0_REG_lrs1_rtype, soc2.core.iregister_read.rrd_uops_0_REG_lrs2_rtype) &&
	check_uopc_lrs1_lrs2(soc2.core.iregister_read.rrd_uops_1_REG_uopc, soc2.core.iregister_read.rrd_uops_1_REG_lrs1_rtype, soc2.core.iregister_read.rrd_uops_1_REG_lrs2_rtype) &&
	check_uopc_lrs1_lrs2(soc2.core.iregister_read.rrd_uops_2_REG_uopc, soc2.core.iregister_read.rrd_uops_2_REG_lrs1_rtype, soc2.core.iregister_read.rrd_uops_2_REG_lrs2_rtype) &&
	check_fp_uopc_lrs1_lrs2(soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_uopc, soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_lrs1_rtype, soc2.core.fp_pipeline.fregister_read.rrd_uops_0_REG_lrs2_rtype);
	
	wire rrd_op_sel_2;
	assign rrd_op_sel_2 =
		check_uopc_op_sel(soc2.core.iregister_read.rrd_uops_1_REG_uopc, soc2.core.iregister_read.rrd_uops_1_REG_ctrl_op1_sel, soc2.core.iregister_read.rrd_uops_1_REG_ctrl_op2_sel) &&
		check_uopc_op_sel(soc2.core.iregister_read.rrd_uops_2_REG_uopc, soc2.core.iregister_read.rrd_uops_2_REG_ctrl_op1_sel, soc2.core.iregister_read.rrd_uops_2_REG_ctrl_op2_sel);
	
	wire csr_alu_req_uopc_2;
	assign csr_alu_req_uopc_2 = !soc2.core.csr_exe_unit.alu.io_req_valid || check_csr_alu_uopc(soc2.core.csr_exe_unit.alu.io_req_bits_uop_uopc);  
	
	wire csr_div_req_uopc_2;
	assign csr_div_req_uopc_2 = !soc2.core.csr_exe_unit.div.io_req_valid || check_csr_div_uopc(soc2.core.csr_exe_unit.div.io_req_bits_uop_uopc);
	
	wire jmp_unit_alu_req_uopc_2;
	assign jmp_unit_alu_req_uopc_2 = !soc2.core.jmp_unit.alu.io_req_valid || check_jmp_unit_alu_uopc(soc2.core.jmp_unit.alu.io_req_bits_uop_uopc);
	
	wire jmp_unit_ifpu_req_uopc_2;
	assign jmp_unit_ifpu_req_uopc_2 = !soc2.core.jmp_unit.ifpu.io_req_valid || check_jmp_unit_ifpu_uopc(soc2.core.jmp_unit.ifpu.io_req_bits_uop_uopc);
	
	wire dmem_resp_equals_s2_type_2;
	assign dmem_resp_equals_s2_type_2 = soc2.lsu.io_dmem_resp_0_valid && soc2.dcache.cache_resp_0_valid ? soc2.dcache.s2_type == 3'h4 || soc2.dcache.s2_type == 3'h0 : 1'b1;
	
	wire s2_hella_matching_s2_type_2;
	assign s2_hella_matching_s2_type_2 = soc2.dcache.s2_valid_REG && soc2.dcache.s2_req_0_is_hella ? soc2.dcache.s2_type == 3'h4 : 1'b1;
	
	wire will_fire_sfence_not_speculative_2;
	assign will_fire_sfence_not_speculative_2 = soc2.lsu.will_fire_sfence_0_will_fire ? soc2.lsu.io_core_exe_0_req_bits_uop_br_mask == 12'h0 : 1'b1;
	
	wire store_req_not_committed_2;
	assign store_req_not_committed_2 = soc2.lsu.io_core_exe_0_req_valid && soc2.lsu.io_core_exe_0_req_bits_uop_uses_stq ? !stq_committed_2[soc2.lsu.io_core_exe_0_req_bits_uop_stq_idx] : 1'b1;
	
	wire hella_not_using_ldq_stq_2;
	assign hella_not_using_ldq_stq_2 = soc2.lsu.io_dmem_resp_0_bits_is_hella ? !soc2.lsu.io_dmem_resp_0_bits_uop_uses_ldq && !soc2.lsu.io_dmem_resp_0_bits_uop_uses_stq : 1'b1;
	
	wire s2_amo_nonspeculative_2;
	assign s2_amo_nonspeculative_2 = soc2.dcache.s2_valid_REG && soc2.dcache.s2_req_0_uop_is_amo ? soc2.dcache.s2_req_0_uop_br_mask == 12'h0 : 1'b1;
	
	wire committed_store_not_being_tainted_2;
	assign committed_store_not_being_tainted_2 =
		//GEN signals can be found by searching for io_core_exe_0_req_valid & io_core_exe_0_req_bits_uop_uses_stq & io_core_exe_0_req_bits_uop_taint ? _GEN_37623 : _GEN_37485; // @[lsu.scala 1580:89]
		(stq_valids_2[0] && stq_committed_2[0] ? !soc2.lsu._GEN_37477 : 1'b1) &&
		(stq_valids_2[1] && stq_committed_2[1] ? !soc2.lsu._GEN_37478 : 1'b1) &&
		(stq_valids_2[2] && stq_committed_2[2] ? !soc2.lsu._GEN_37479 : 1'b1) &&
		(stq_valids_2[3] && stq_committed_2[3] ? !soc2.lsu._GEN_37480 : 1'b1) &&
		(stq_valids_2[4] && stq_committed_2[4] ? !soc2.lsu._GEN_37481 : 1'b1) &&
		(stq_valids_2[5] && stq_committed_2[5] ? !soc2.lsu._GEN_37482 : 1'b1) &&
		(stq_valids_2[6] && stq_committed_2[6] ? !soc2.lsu._GEN_37483 : 1'b1) &&
		(stq_valids_2[7] && stq_committed_2[7] ? !soc2.lsu._GEN_37484 : 1'b1) &&
		(stq_valids_2[8] && stq_committed_2[8] ? !soc2.lsu._GEN_37485 : 1'b1) &&
		(stq_valids_2[9] && stq_committed_2[9] ? !soc2.lsu._GEN_37486 : 1'b1) &&
		(stq_valids_2[10] && stq_committed_2[10] ? !soc2.lsu._GEN_37487 : 1'b1) &&
		(stq_valids_2[11] && stq_committed_2[11] ? !soc2.lsu._GEN_37488 : 1'b1) &&
		(stq_valids_2[12] && stq_committed_2[12] ? !soc2.lsu._GEN_37489 : 1'b1) &&
		(stq_valids_2[13] && stq_committed_2[13] ? !soc2.lsu._GEN_37490 : 1'b1) &&
		(stq_valids_2[14] && stq_committed_2[14] ? !soc2.lsu._GEN_37491 : 1'b1) &&
		(stq_valids_2[15] && stq_committed_2[15] ? !soc2.lsu._GEN_37492 : 1'b1);
		
	wire exe_reg_0_sfence_not_speculative_2;
	assign exe_reg_0_sfence_not_speculative_2 = soc2.core.iregister_read.exe_reg_valids_0 && soc2.core.iregister_read.exe_reg_uops_0_mem_cmd == 5'h14 ? soc2.core.iregister_read.exe_reg_uops_0_br_mask == 12'h0 : 1'b1; 
	
	wire rrd_no_rocc_2;
	assign rrd_no_rocc_2 =
	(soc2.core.iregister_read.rrd_uops_0_REG_uopc != 7'h6c) && (soc2.core.iregister_read.rrd_uops_1_REG_uopc != 7'h6c) && (soc2.core.iregister_read.rrd_uops_2_REG_uopc != 7'h6c);
	
	wire dmem_req_amo_2;
	assign dmem_req_amo_2 = soc2.lsu.io_dmem_req_bits_0_valid && soc2.lsu.io_dmem_req_bits_0_bits_uop_is_amo? soc2.lsu.io_dmem_req_bits_0_bits_uop_br_mask == 12'h0 : 1'b1;
	
	wire fpu_req_uopc_2;
	assign fpu_req_uopc_2 = !soc2.core.fp_pipeline.fpiu_unit.fpu.io_req_valid || check_fpu_uopc(soc2.core.fp_pipeline.fpiu_unit.fpu.io_req_bits_uop_uopc);
	
	wire fdivsqrt_req_uopc_2;
	assign fdivsqrt_req_uopc_2 = !soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.io_req_valid || check_fdivsqrt_uopc(soc2.core.fp_pipeline.fpiu_unit.fdivsqrt.io_req_bits_uop_uopc);
	
	wire fp_sdq_req_uopc_2;
	assign fp_sdq_req_uopc_2 = !soc2.core.fp_pipeline.fpiu_unit.fp_sdq.io_enq_valid || soc2.core.fp_pipeline.fpiu_unit.fp_sdq.io_enq_bits_uop_uopc == 7'h2;
	
	wire br_jal_jalr_consistent_uopc_2;
	assign br_jal_jalr_consistent_uopc_2 =
	(soc2.core.iregister_read.exe_reg_uops_1_is_br
	?
		soc2.core.iregister_read.exe_reg_uops_1_uopc == 7'h18 || soc2.core.iregister_read.exe_reg_uops_1_uopc == 7'h19 || soc2.core.iregister_read.exe_reg_uops_1_uopc == 7'h1a ||
		soc2.core.iregister_read.exe_reg_uops_1_uopc == 7'h1b || soc2.core.iregister_read.exe_reg_uops_1_uopc == 7'h1c || soc2.core.iregister_read.exe_reg_uops_1_uopc == 7'h1d
	: 1'b1) &&
	(soc2.core.iregister_read.exe_reg_uops_1_is_jal ? soc2.core.iregister_read.exe_reg_uops_1_uopc == 7'h25 : 1'b1) &&
	(soc2.core.iregister_read.exe_reg_uops_1_is_jalr ? soc2.core.iregister_read.exe_reg_uops_1_uopc == 7'h26 : 1'b1) &&
	(soc2.core.iregister_read.exe_reg_uops_2_is_br
	?
		soc2.core.iregister_read.exe_reg_uops_2_uopc == 7'h18 || soc2.core.iregister_read.exe_reg_uops_2_uopc == 7'h19 || soc2.core.iregister_read.exe_reg_uops_2_uopc == 7'h1a ||
		soc2.core.iregister_read.exe_reg_uops_2_uopc == 7'h1b || soc2.core.iregister_read.exe_reg_uops_2_uopc == 7'h1c || soc2.core.iregister_read.exe_reg_uops_2_uopc == 7'h1d
	: 1'b1) &&
	(soc2.core.iregister_read.exe_reg_uops_2_is_jal ? soc2.core.iregister_read.exe_reg_uops_2_uopc == 7'h25 : 1'b1) &&
	(soc2.core.iregister_read.exe_reg_uops_2_is_jalr ? soc2.core.iregister_read.exe_reg_uops_2_uopc == 7'h26 : 1'b1);

	//br_type and uopc consistent
	wire br_type_consistent_2;
	assign br_type_consistent_2 =
		(soc2.core.iregister_read.exe_reg_uops_1_ctrl_br_type == 4'h8 ? soc2.core.iregister_read.exe_reg_uops_1_uopc == 7'h26 : 1'b1) &&
    		(soc2.core.iregister_read.exe_reg_uops_2_ctrl_br_type == 4'h8 ? soc2.core.iregister_read.exe_reg_uops_2_uopc == 7'h26 : 1'b1);
    	    
    	wire sfence_at_head_2;
    	assign sfence_at_head_2 =
    		soc2.core.mem_units_0.maddrcalc.io_resp_bits_sfence_valid ? soc2.core.mem_units_0.maddrcalc.io_resp_bits_uop_rob_idx == soc2.core.rob.io_rob_head_idx : 1'b1;
	
	//wire ifpu_valids_consistent_2;
	//assign ifpu_valids_consistent_2 = soc2.core.jmp_unit.ifpu.ifpu.io_out_v ? soc2.core.jmp_unit.ifpu.r_valids_1 : 1'b1;
	
	wire fp_exe_reg_yrot;
	assign fp_exe_reg_yrot =
		(soc1.core.fp_pipeline.fregister_read.exe_reg_rs1_data_0 != soc2.core.fp_pipeline.fregister_read.exe_reg_rs1_data_0 ||
		soc1.core.fp_pipeline.fregister_read.exe_reg_rs2_data_0 != soc2.core.fp_pipeline.fregister_read.exe_reg_rs2_data_0 ||
		soc1.core.fp_pipeline.fregister_read.exe_reg_rs3_data_0 != soc2.core.fp_pipeline.fregister_read.exe_reg_rs3_data_0) 
		? 
			ROBisOlder(soc1.core.rob.io_rob_pnr_idx, soc1.core.fp_pipeline.fregister_read.exe_reg_yrot_0, soc1.core.rob.io_rob_head_idx) &&
			ROBisOlder(soc2.core.rob.io_rob_pnr_idx, soc2.core.fp_pipeline.fregister_read.exe_reg_yrot_0, soc2.core.rob.io_rob_head_idx) 
		: 1'b1;
		
	wire int_exe_reg_yrot;
	assign int_exe_reg_yrot =
		(
			(soc1.core.iregister_read.exe_reg_rs1_data_0 != soc2.core.iregister_read.exe_reg_rs1_data_0 ||
			soc1.core.iregister_read.exe_reg_rs2_data_0 != soc2.core.iregister_read.exe_reg_rs2_data_0) 
			? 
				ROBisOlder(soc1.core.rob.io_rob_pnr_idx, soc1.core.iregister_read.exe_reg_yrot_0, soc1.core.rob.io_rob_head_idx) &&
				ROBisOlder(soc2.core.rob.io_rob_pnr_idx, soc2.core.iregister_read.exe_reg_yrot_0, soc2.core.rob.io_rob_head_idx) 
			: 1'b1
		) &&
		(
			(soc1.core.iregister_read.exe_reg_rs1_data_1 != soc2.core.iregister_read.exe_reg_rs1_data_1 ||
			soc1.core.iregister_read.exe_reg_rs2_data_1 != soc2.core.iregister_read.exe_reg_rs2_data_1) 
			? 
				ROBisOlder(soc1.core.rob.io_rob_pnr_idx, soc1.core.iregister_read.exe_reg_yrot_1, soc1.core.rob.io_rob_head_idx) &&
				ROBisOlder(soc2.core.rob.io_rob_pnr_idx, soc2.core.iregister_read.exe_reg_yrot_1, soc2.core.rob.io_rob_head_idx) 
			: 1'b1
		) &&
		(
			(soc1.core.iregister_read.exe_reg_rs1_data_2 != soc2.core.iregister_read.exe_reg_rs1_data_2 ||
			soc1.core.iregister_read.exe_reg_rs2_data_2 != soc2.core.iregister_read.exe_reg_rs2_data_2) 
			? 
				ROBisOlder(soc1.core.rob.io_rob_pnr_idx, soc1.core.iregister_read.exe_reg_yrot_2, soc1.core.rob.io_rob_head_idx) &&
				ROBisOlder(soc2.core.rob.io_rob_pnr_idx, soc2.core.iregister_read.exe_reg_yrot_2, soc2.core.rob.io_rob_head_idx) 
			: 1'b1
		);
	
	wire dmem_resp_uncommittable;
	assign dmem_resp_uncommittable = 
	soc1.lsu.io_dmem_resp_0_valid && soc1.lsu.io_dmem_resp_0_bits_uop_uses_ldq && soc2.lsu.io_dmem_resp_0_valid && soc2.lsu.io_dmem_resp_0_bits_uop_uses_ldq &&
	(soc1.lsu.io_dmem_resp_0_bits_uop_ldq_idx == soc2.lsu.io_dmem_resp_0_bits_uop_ldq_idx) &&
	(soc1.lsu.io_dmem_resp_0_bits_data != soc2.lsu.io_dmem_resp_0_bits_data)
	?
		!ROBisOlder(ldq_rob_idx_1,root_id,soc1.core.rob.io_rob_head_idx) && 
		!ROBisOlder(ldq_rob_idx_2,root_id,soc2.core.rob.io_rob_head_idx)
	:
		1'b1;
		
	wire ptw_not_accessing_secret;
	assign ptw_not_accessing_secret =
   		(soc1.dcache.s2_valid_REG && soc1.dcache.s2_req_0_is_hella ? soc1.dcache.s2_req_0_addr[31:12] != 20'h8abcd : 1'b1) && 
   		(soc2.dcache.s2_valid_REG && soc2.dcache.s2_req_0_is_hella ? soc2.dcache.s2_req_0_addr[31:12] != 20'h8abcd : 1'b1); 
   		
   	wire ifpu_out_uncommittable;
   	assign ifpu_out_uncommittable =
   		soc1.core.jmp_unit.ifpu.r_uops_1_rob_idx == soc2.core.jmp_unit.ifpu.r_uops_1_rob_idx &&
   		soc1.core.jmp_unit.ifpu.ifpu.io_out_b_exc != soc2.core.jmp_unit.ifpu.ifpu.io_out_b_exc
   		?
   			!isRobIdCommitable(soc1.core.rob.rob_head, root_id, soc1.core.jmp_unit.ifpu.r_uops_1_rob_idx) &&
   			!isRobIdCommitable(soc2.core.rob.rob_head, root_id, soc2.core.jmp_unit.ifpu.r_uops_1_rob_idx)
		:
			1'b1;
			
	wire rob_fflags_uncommittable;
	assign rob_fflags_uncommittable =
		(soc1.core.rob.rob_fflags[0] != soc2.core.rob.rob_fflags[0] ? ROBisOlder(root_id,6'h0,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h0,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h0 && soc2.core.rob.io_rob_head_idx != 6'h0 && (rob_branch_masks_1[6'h0] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h0] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[1] != soc2.core.rob.rob_fflags[1] ? ROBisOlder(root_id,6'h2,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h2,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h2 && soc2.core.rob.io_rob_head_idx != 6'h2 && (rob_branch_masks_1[6'h2] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h2] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[2] != soc2.core.rob.rob_fflags[2] ? ROBisOlder(root_id,6'h4,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h4,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h4 && soc2.core.rob.io_rob_head_idx != 6'h4 && (rob_branch_masks_1[6'h4] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h4] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[3] != soc2.core.rob.rob_fflags[3] ? ROBisOlder(root_id,6'h6,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h6,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h6 && soc2.core.rob.io_rob_head_idx != 6'h6 && (rob_branch_masks_1[6'h6] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h6] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[4] != soc2.core.rob.rob_fflags[4] ? ROBisOlder(root_id,6'h8,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h8,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h8 && soc2.core.rob.io_rob_head_idx != 6'h8 && (rob_branch_masks_1[6'h8] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h8] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[5] != soc2.core.rob.rob_fflags[5] ? ROBisOlder(root_id,6'ha,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'ha,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'ha && soc2.core.rob.io_rob_head_idx != 6'ha && (rob_branch_masks_1[6'ha] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'ha] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[6] != soc2.core.rob.rob_fflags[6] ? ROBisOlder(root_id,6'hc,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'hc,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'hc && soc2.core.rob.io_rob_head_idx != 6'hc && (rob_branch_masks_1[6'hc] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'hc] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[7] != soc2.core.rob.rob_fflags[7] ? ROBisOlder(root_id,6'he,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'he,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'he && soc2.core.rob.io_rob_head_idx != 6'he && (rob_branch_masks_1[6'he] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'he] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[8] != soc2.core.rob.rob_fflags[8] ? ROBisOlder(root_id,6'h10,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h10,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h10 && soc2.core.rob.io_rob_head_idx != 6'h10 && (rob_branch_masks_1[6'h10] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h10] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[9] != soc2.core.rob.rob_fflags[9] ? ROBisOlder(root_id,6'h12,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h12,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h12 && soc2.core.rob.io_rob_head_idx != 6'h12 && (rob_branch_masks_1[6'h12] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h12] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[10] != soc2.core.rob.rob_fflags[10] ? ROBisOlder(root_id,6'h14,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h14,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h14 && soc2.core.rob.io_rob_head_idx != 6'h14 && (rob_branch_masks_1[6'h14] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h14] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[11] != soc2.core.rob.rob_fflags[11] ? ROBisOlder(root_id,6'h16,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h16,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h16 && soc2.core.rob.io_rob_head_idx != 6'h16 && (rob_branch_masks_1[6'h16] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h16] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[12] != soc2.core.rob.rob_fflags[12] ? ROBisOlder(root_id,6'h18,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h18,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h18 && soc2.core.rob.io_rob_head_idx != 6'h18 && (rob_branch_masks_1[6'h18] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h18] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[13] != soc2.core.rob.rob_fflags[13] ? ROBisOlder(root_id,6'h1a,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h1a,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h1a && soc2.core.rob.io_rob_head_idx != 6'h1a && (rob_branch_masks_1[6'h1a] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h1a] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[14] != soc2.core.rob.rob_fflags[14] ? ROBisOlder(root_id,6'h1c,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h1c,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h1c && soc2.core.rob.io_rob_head_idx != 6'h1c && (rob_branch_masks_1[6'h1c] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h1c] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[15] != soc2.core.rob.rob_fflags[15] ? ROBisOlder(root_id,6'h1e,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h1e,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h1e && soc2.core.rob.io_rob_head_idx != 6'h1e && (rob_branch_masks_1[6'h1e] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h1e] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[16] != soc2.core.rob.rob_fflags[16] ? ROBisOlder(root_id,6'h20,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h20,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h20 && soc2.core.rob.io_rob_head_idx != 6'h20 && (rob_branch_masks_1[6'h20] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h20] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[17] != soc2.core.rob.rob_fflags[17] ? ROBisOlder(root_id,6'h22,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h22,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h22 && soc2.core.rob.io_rob_head_idx != 6'h22 && (rob_branch_masks_1[6'h22] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h22] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[18] != soc2.core.rob.rob_fflags[18] ? ROBisOlder(root_id,6'h24,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h24,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h24 && soc2.core.rob.io_rob_head_idx != 6'h24 && (rob_branch_masks_1[6'h24] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h24] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[19] != soc2.core.rob.rob_fflags[19] ? ROBisOlder(root_id,6'h26,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h26,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h26 && soc2.core.rob.io_rob_head_idx != 6'h26 && (rob_branch_masks_1[6'h26] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h26] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[20] != soc2.core.rob.rob_fflags[20] ? ROBisOlder(root_id,6'h28,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h28,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h28 && soc2.core.rob.io_rob_head_idx != 6'h28 && (rob_branch_masks_1[6'h28] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h28] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[21] != soc2.core.rob.rob_fflags[21] ? ROBisOlder(root_id,6'h2a,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h2a,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h2a && soc2.core.rob.io_rob_head_idx != 6'h2a && (rob_branch_masks_1[6'h2a] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h2a] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[22] != soc2.core.rob.rob_fflags[22] ? ROBisOlder(root_id,6'h2c,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h2c,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h2c && soc2.core.rob.io_rob_head_idx != 6'h2c && (rob_branch_masks_1[6'h2c] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h2c] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[23] != soc2.core.rob.rob_fflags[23] ? ROBisOlder(root_id,6'h2e,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h2e,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h2e && soc2.core.rob.io_rob_head_idx != 6'h2e && (rob_branch_masks_1[6'h2e] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h2e] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[24] != soc2.core.rob.rob_fflags[24] ? ROBisOlder(root_id,6'h30,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h30,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h30 && soc2.core.rob.io_rob_head_idx != 6'h30 && (rob_branch_masks_1[6'h30] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h30] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[25] != soc2.core.rob.rob_fflags[25] ? ROBisOlder(root_id,6'h32,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h32,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h32 && soc2.core.rob.io_rob_head_idx != 6'h32 && (rob_branch_masks_1[6'h32] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h32] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[26] != soc2.core.rob.rob_fflags[26] ? ROBisOlder(root_id,6'h34,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h34,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h34 && soc2.core.rob.io_rob_head_idx != 6'h34 && (rob_branch_masks_1[6'h34] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h34] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[27] != soc2.core.rob.rob_fflags[27] ? ROBisOlder(root_id,6'h36,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h36,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h36 && soc2.core.rob.io_rob_head_idx != 6'h36 && (rob_branch_masks_1[6'h36] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h36] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[28] != soc2.core.rob.rob_fflags[28] ? ROBisOlder(root_id,6'h38,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h38,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h38 && soc2.core.rob.io_rob_head_idx != 6'h38 && (rob_branch_masks_1[6'h38] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h38] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[29] != soc2.core.rob.rob_fflags[29] ? ROBisOlder(root_id,6'h3a,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h3a,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h3a && soc2.core.rob.io_rob_head_idx != 6'h3a && (rob_branch_masks_1[6'h3a] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h3a] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[30] != soc2.core.rob.rob_fflags[30] ? ROBisOlder(root_id,6'h3c,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h3c,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h3c && soc2.core.rob.io_rob_head_idx != 6'h3c && (rob_branch_masks_1[6'h3c] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h3c] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags[31] != soc2.core.rob.rob_fflags[31] ? ROBisOlder(root_id,6'h3e,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h3e,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h3e && soc2.core.rob.io_rob_head_idx != 6'h3e && (rob_branch_masks_1[6'h3e] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h3e] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[0] != soc2.core.rob.rob_fflags_1[0] ? ROBisOlder(root_id,6'h1,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h1,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h1 && soc2.core.rob.io_rob_head_idx != 6'h1 && (rob_branch_masks_1[6'h1] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h1] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[1] != soc2.core.rob.rob_fflags_1[1] ? ROBisOlder(root_id,6'h3,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h3,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h3 && soc2.core.rob.io_rob_head_idx != 6'h3 && (rob_branch_masks_1[6'h3] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h3] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[2] != soc2.core.rob.rob_fflags_1[2] ? ROBisOlder(root_id,6'h5,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h5,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h5 && soc2.core.rob.io_rob_head_idx != 6'h5 && (rob_branch_masks_1[6'h5] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h5] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[3] != soc2.core.rob.rob_fflags_1[3] ? ROBisOlder(root_id,6'h7,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h7,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h7 && soc2.core.rob.io_rob_head_idx != 6'h7 && (rob_branch_masks_1[6'h7] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h7] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[4] != soc2.core.rob.rob_fflags_1[4] ? ROBisOlder(root_id,6'h9,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h9,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h9 && soc2.core.rob.io_rob_head_idx != 6'h9 && (rob_branch_masks_1[6'h9] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h9] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[5] != soc2.core.rob.rob_fflags_1[5] ? ROBisOlder(root_id,6'hb,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'hb,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'hb && soc2.core.rob.io_rob_head_idx != 6'hb && (rob_branch_masks_1[6'hb] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'hb] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[6] != soc2.core.rob.rob_fflags_1[6] ? ROBisOlder(root_id,6'hd,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'hd,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'hd && soc2.core.rob.io_rob_head_idx != 6'hd && (rob_branch_masks_1[6'hd] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'hd] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[7] != soc2.core.rob.rob_fflags_1[7] ? ROBisOlder(root_id,6'hf,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'hf,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'hf && soc2.core.rob.io_rob_head_idx != 6'hf && (rob_branch_masks_1[6'hf] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'hf] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[8] != soc2.core.rob.rob_fflags_1[8] ? ROBisOlder(root_id,6'h11,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h11,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h11 && soc2.core.rob.io_rob_head_idx != 6'h11 && (rob_branch_masks_1[6'h11] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h11] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[9] != soc2.core.rob.rob_fflags_1[9] ? ROBisOlder(root_id,6'h13,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h13,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h13 && soc2.core.rob.io_rob_head_idx != 6'h13 && (rob_branch_masks_1[6'h13] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h13] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[10] != soc2.core.rob.rob_fflags_1[10] ? ROBisOlder(root_id,6'h15,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h15,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h15 && soc2.core.rob.io_rob_head_idx != 6'h15 && (rob_branch_masks_1[6'h15] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h15] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[11] != soc2.core.rob.rob_fflags_1[11] ? ROBisOlder(root_id,6'h17,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h17,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h17 && soc2.core.rob.io_rob_head_idx != 6'h17 && (rob_branch_masks_1[6'h17] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h17] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[12] != soc2.core.rob.rob_fflags_1[12] ? ROBisOlder(root_id,6'h19,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h19,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h19 && soc2.core.rob.io_rob_head_idx != 6'h19 && (rob_branch_masks_1[6'h19] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h19] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[13] != soc2.core.rob.rob_fflags_1[13] ? ROBisOlder(root_id,6'h1b,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h1b,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h1b && soc2.core.rob.io_rob_head_idx != 6'h1b && (rob_branch_masks_1[6'h1b] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h1b] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[14] != soc2.core.rob.rob_fflags_1[14] ? ROBisOlder(root_id,6'h1d,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h1d,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h1d && soc2.core.rob.io_rob_head_idx != 6'h1d && (rob_branch_masks_1[6'h1d] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h1d] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[15] != soc2.core.rob.rob_fflags_1[15] ? ROBisOlder(root_id,6'h1f,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h1f,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h1f && soc2.core.rob.io_rob_head_idx != 6'h1f && (rob_branch_masks_1[6'h1f] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h1f] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[16] != soc2.core.rob.rob_fflags_1[16] ? ROBisOlder(root_id,6'h21,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h21,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h21 && soc2.core.rob.io_rob_head_idx != 6'h21 && (rob_branch_masks_1[6'h21] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h21] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[17] != soc2.core.rob.rob_fflags_1[17] ? ROBisOlder(root_id,6'h23,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h23,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h23 && soc2.core.rob.io_rob_head_idx != 6'h23 && (rob_branch_masks_1[6'h23] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h23] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[18] != soc2.core.rob.rob_fflags_1[18] ? ROBisOlder(root_id,6'h25,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h25,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h25 && soc2.core.rob.io_rob_head_idx != 6'h25 && (rob_branch_masks_1[6'h25] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h25] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[19] != soc2.core.rob.rob_fflags_1[19] ? ROBisOlder(root_id,6'h27,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h27,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h27 && soc2.core.rob.io_rob_head_idx != 6'h27 && (rob_branch_masks_1[6'h27] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h27] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[20] != soc2.core.rob.rob_fflags_1[20] ? ROBisOlder(root_id,6'h29,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h29,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h29 && soc2.core.rob.io_rob_head_idx != 6'h29 && (rob_branch_masks_1[6'h29] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h29] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[21] != soc2.core.rob.rob_fflags_1[21] ? ROBisOlder(root_id,6'h2b,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h2b,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h2b && soc2.core.rob.io_rob_head_idx != 6'h2b && (rob_branch_masks_1[6'h2b] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h2b] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[22] != soc2.core.rob.rob_fflags_1[22] ? ROBisOlder(root_id,6'h2d,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h2d,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h2d && soc2.core.rob.io_rob_head_idx != 6'h2d && (rob_branch_masks_1[6'h2d] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h2d] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[23] != soc2.core.rob.rob_fflags_1[23] ? ROBisOlder(root_id,6'h2f,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h2f,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h2f && soc2.core.rob.io_rob_head_idx != 6'h2f && (rob_branch_masks_1[6'h2f] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h2f] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[24] != soc2.core.rob.rob_fflags_1[24] ? ROBisOlder(root_id,6'h31,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h31,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h31 && soc2.core.rob.io_rob_head_idx != 6'h31 && (rob_branch_masks_1[6'h31] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h31] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[25] != soc2.core.rob.rob_fflags_1[25] ? ROBisOlder(root_id,6'h33,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h33,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h33 && soc2.core.rob.io_rob_head_idx != 6'h33 && (rob_branch_masks_1[6'h33] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h33] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[26] != soc2.core.rob.rob_fflags_1[26] ? ROBisOlder(root_id,6'h35,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h35,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h35 && soc2.core.rob.io_rob_head_idx != 6'h35 && (rob_branch_masks_1[6'h35] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h35] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[27] != soc2.core.rob.rob_fflags_1[27] ? ROBisOlder(root_id,6'h37,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h37,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h37 && soc2.core.rob.io_rob_head_idx != 6'h37 && (rob_branch_masks_1[6'h37] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h37] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[28] != soc2.core.rob.rob_fflags_1[28] ? ROBisOlder(root_id,6'h39,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h39,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h39 && soc2.core.rob.io_rob_head_idx != 6'h39 && (rob_branch_masks_1[6'h39] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h39] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[29] != soc2.core.rob.rob_fflags_1[29] ? ROBisOlder(root_id,6'h3b,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h3b,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h3b && soc2.core.rob.io_rob_head_idx != 6'h3b && (rob_branch_masks_1[6'h3b] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h3b] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[30] != soc2.core.rob.rob_fflags_1[30] ? ROBisOlder(root_id,6'h3d,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h3d,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h3d && soc2.core.rob.io_rob_head_idx != 6'h3d && (rob_branch_masks_1[6'h3d] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h3d] & root_br_mask) != 12'h0 : 1'b1) &&
		(soc1.core.rob.rob_fflags_1[31] != soc2.core.rob.rob_fflags_1[31] ? ROBisOlder(root_id,6'h3f,soc1.core.rob.io_rob_head_idx) && ROBisOlder(root_id,6'h3f,soc2.core.rob.io_rob_head_idx) && soc1.core.rob.io_rob_head_idx != 6'h3f && soc2.core.rob.io_rob_head_idx != 6'h3f && (rob_branch_masks_1[6'h3f] & root_br_mask) != 12'h0 && (rob_branch_masks_2[6'h3f] & root_br_mask) != 12'h0 : 1'b1);	

	//arrays for symbolic proof commitment
	wire ROB_commit_array_1 [1:0];
	assign ROB_commit_array_1[0] = soc1.core.rob.io_commit_valids_0;
	assign ROB_commit_array_1[1] = soc1.core.rob.io_commit_valids_1;
	
	wire ROB_commit_array_2 [1:0];
	assign ROB_commit_array_2[0] = soc2.core.rob.io_commit_valids_0;
	assign ROB_commit_array_2[1] = soc2.core.rob.io_commit_valids_1;
	

endmodule

	// This is based on the assumption that the ability of attacker to measure
	// time is synchronized with instruction commit
	// in case of RISC-V csr timers: csr reads are synchronizing instructions
	// in case of external timers: signaling the outside world should never be
	// done speculatively
	// if timer reading is not synchronized: the upec L-Alert definition becomes
	// even more simple, i.e., every physical register can be considered
	// architectural, but it becomes extremely hard to have a secure variant
	// it may not also make sense to allow SW to measure time in such a fine
	// grained manner
